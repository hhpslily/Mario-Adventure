module pixel_gen(
	input clk,
    input rst,
	input valid,
	input [2:0] state,
    input [9:0] h_cnt,
    input [9:0] v_cnt,
    input [9:0] x, 
    input [11:0] pixel,
	
	output reg die,
	output reg [2:0] LED,
    output reg [3:0] vgaRed,
    output reg [3:0] vgaGreen,
    output reg [3:0] vgaBlue,
	output reg [11:0] point
   );
	
	reg point1,point2,point3,point4,point5;
	reg [1:0] life;
	reg [9:0] bagel1_x, bagel1_y, bagel2_x, bagel2_y, bagel3_x, bagel3_y, bagel4_x, bagel4_y, bagel5_x, bagel5_y, 
	          branch1_x, branch1_y,branch2_x, branch2_y,branch3_x, branch3_y,branch4_x, branch4_y,branch5_x, branch5_y;
    reg [30:0] num;
    wire [30:0] next_num;
    always @(posedge clk) begin
          num <= next_num;
    end
    assign next_num = num + 1'b1;
    always @ (posedge clk or posedge rst) begin
        if(rst) begin
            bagel1_x <= 29;
            bagel1_y <= 0;
            bagel2_x <= 165;
            bagel2_y <= -473;
            bagel3_x <= 301;
            bagel3_y <= -328;
            bagel4_x <= 437;
            bagel4_y <= -183;
            bagel5_x <= 573;
            bagel5_y <= -294;
            branch1_x <= 29;
            branch1_y <= -597;
            branch2_x <= 165;
            branch2_y <= -177;
            branch3_x <= 301;
            branch3_y <= -666;
            branch4_x <= 437;
            branch4_y <= -920;
            branch5_x <= 573;
            branch5_y <= -777;
			point1<= 0;
			point2<= 0;
			point3<= 0;
			point4<= 0;
			point5<= 0;
			life<=3;
			die<=0;
        end else begin
			if(bagel1_y==324 && x==bagel1_x-29)begin
				bagel1_y <= 0;
				point1<=1;				
			end else if(branch1_y==322 && x==branch1_x-29) begin
				branch1_y <= -597;
				point1<=0;
				if(life>=1)
					life<=life-1;
				else
					die<=1;
			end else begin
				bagel1_y <= (state!=3'b011)?bagel1_y+1:bagel1_y;
				branch1_y <= (state!=3'b011)?branch1_y+1:branch1_y;
				point1<=0;
			end
            
			if(bagel2_y==324 && x==bagel2_x-29)begin
				bagel2_y <= -473;
				point2<=1;
            end else if(branch2_y==322 && x==branch2_x-29) begin
				branch2_y <= -177;
				point2<=0;
				if(life>=1)
					life<=life-1;
				else
					die<=1;
			end else begin
      			bagel2_y <= (state!=3'b011)?bagel2_y+1:bagel2_y;
				branch2_y <= (state!=3'b011)?branch2_y+1:branch2_y;
      			point2<=0;
      		end
            
			if(bagel3_y==324 && x==bagel3_x-29)begin
				bagel3_y <= -328;
				point3<=1;
            end else if(branch3_y==322 && x==branch3_x-29) begin
				branch3_y <= -666;
				point3<=0;
				if(life>=1)
					life<=life-1;
				else
					die<=1;
			end else begin
            	bagel3_y <= (state!=3'b011)?bagel3_y+1:bagel3_y;
				branch3_y <= (state!=3'b011)?branch3_y+1:branch3_y;
            	point3<=0;
            end
            
			if(bagel4_y==324 && x==bagel4_x-29)begin
				bagel4_y <= -183;
				point4<=1;
            end else if(branch4_y==322 && x==branch4_x-29) begin
				branch4_y <= -929;
				point4<=0;
				if(life>=1)
					life<=life-1;
				else
					die<=1;
			end else begin
            	bagel4_y <= (state!=3'b011)?bagel4_y+1:bagel4_y;
				branch4_y <= (state!=3'b011)?branch4_y+1:branch4_y;
            	point4<=0;
            end
            
			if(bagel5_y==324 && x==bagel5_x-29)begin
				bagel5_y <= -294;
				point5<=1;
            end else if(branch5_y==322 && x==branch5_x-29) begin
				branch5_y <= -777;
				point5<=0;
				if(life>=1)
					life<=life-1;
				else
					die<=1;
			end else begin
            	bagel5_y <= (state!=3'b011)?bagel5_y+1:bagel5_y;
				branch5_y <= (state!=3'b011)?branch5_y+1:branch5_y;
            	point5<=0;
            end
        end
    end
	
	always @(posedge clk) begin
        if(rst) begin
			point<=12'b0;
        end else begin
			point<=(state==3'b001 && point<626)?point1+point2+point3+point4+point5+point:point;
        end
    end
	
	always @* begin	
        if(rst) LED=3'b000;
        else if(life==3) LED=3'b111;
        else if(life==2) LED=3'b011;
        else if(life==1) LED=3'b001;
        else LED=3'b000;
    end
	
	always @(*) begin
		case(state)
			3'b000:begin
				case(num[5])
                                1'b0:begin
                                    if(!valid)
                                        {vgaRed, vgaGreen, vgaBlue} = 12'h0;
                                    else if((((h_cnt >= 80 && h_cnt <= 100) || (h_cnt >= 120 && h_cnt <= 140) || (h_cnt >= 160 && h_cnt <= 180)) && (v_cnt >= 60 && v_cnt <= 200)) || (((h_cnt >= 100 && h_cnt <= 120) || (h_cnt >= 140 && h_cnt <= 160)) && (v_cnt >= 60 && v_cnt <= 80)))
                                        {vgaRed, vgaGreen, vgaBlue} = 12'h39f; // M
                                    else if((((h_cnt >= 200 && h_cnt <= 220) || (h_cnt >= 280 && h_cnt <= 300)) && (v_cnt >= 60 && v_cnt <= 140)) || (((h_cnt >= 220 && h_cnt <= 240) || (h_cnt >= 260 && h_cnt <= 280)) && (v_cnt >= 120 && v_cnt <=140)) || ((h_cnt >= 240 && h_cnt <= 260) && (v_cnt >= 120 && v_cnt <= 220)))
                                         {vgaRed, vgaGreen, vgaBlue} = 12'h0ff; // Y
                                    else if((h_cnt >= 80 && h_cnt <= 100 && v_cnt >= 280 && v_cnt <= 420) || (h_cnt >= 100 && h_cnt <=140 && ((v_cnt >= 280 && v_cnt <= 300) || (v_cnt >= 340 && v_cnt <= 360) || (v_cnt >= 400 && v_cnt <= 420))) ||  (h_cnt >= 140 && h_cnt <= 160 && ((v_cnt >= 300 && v_cnt <= 340) || (v_cnt >= 360 && v_cnt <= 400))))
                                         {vgaRed, vgaGreen, vgaBlue} = 12'h6f6; // B
                                    else if((((h_cnt >= 180 && h_cnt <= 200) || (h_cnt >= 240 && h_cnt <= 260)) && (v_cnt >= 280 && v_cnt <= 420)) || ((h_cnt >= 200 && h_cnt <= 260) && ((v_cnt >= 280 && v_cnt <=300) || (v_cnt >= 340 && v_cnt <=360))))
                                         {vgaRed, vgaGreen, vgaBlue} = 12'hff0; // A              
                                    else if((h_cnt >= 280 && h_cnt <= 300 && v_cnt >= 280 && v_cnt <= 420) || ((h_cnt >= 300 && h_cnt <= 360) && ((v_cnt >= 280 && v_cnt <= 300) || (v_cnt >= 400 && v_cnt <= 420))) || ((h_cnt >= 320 && h_cnt <= 360) && (v_cnt >= 340 && v_cnt <= 360)) || (h_cnt >= 340 && h_cnt <= 360 && v_cnt >= 360 && v_cnt <= 400))
                                         {vgaRed, vgaGreen, vgaBlue} = 12'hf90; // G
                                    else if((h_cnt >= 380 && h_cnt <= 400 && v_cnt >= 280 && v_cnt <= 420) || ((h_cnt >= 400 && h_cnt <= 460) && ((v_cnt >= 280 && v_cnt <= 300) || (v_cnt >= 340 && v_cnt <= 360) || (v_cnt >= 400 && v_cnt <= 420))))
                                         {vgaRed, vgaGreen, vgaBlue} = 12'hf00; // E
                                    else if((h_cnt >= 480 && h_cnt <= 500 && v_cnt >= 280 && v_cnt <= 420) || (h_cnt >= 500 && h_cnt <= 560 && v_cnt >= 400 && v_cnt <= 420))
                                         {vgaRed, vgaGreen, vgaBlue} = 12'hf9c; // L
                                    else if((((h_cnt >= 380 && h_cnt <= 400) || (h_cnt >= 500 && h_cnt <= 520)) && v_cnt >= 100 && v_cnt <= 180) || (h_cnt >= 420 && h_cnt <= 480 && ((v_cnt >= 60 && v_cnt <= 80) || (v_cnt >= 200 && v_cnt <= 220))) || (h_cnt >= 400 && h_cnt <= 420 && v_cnt >= 80 && v_cnt <= 100) || (h_cnt >= 480 && h_cnt <= 500 && v_cnt >= 80 && v_cnt <= 100) || (h_cnt >= 400 && h_cnt <= 420 && v_cnt >= 180 && v_cnt <= 200) || (h_cnt >= 480 && h_cnt <= 500 && v_cnt >= 180 && v_cnt <= 200)) 
                                         {vgaRed, vgaGreen, vgaBlue} = 12'hfff; // bagel(out)
                                    else if((h_cnt >= 420 && h_cnt <= 440 && v_cnt >= 120 && v_cnt <= 160) || (h_cnt >= 460 && h_cnt <= 480 && v_cnt >= 120 && v_cnt <= 160) || (h_cnt >= 440 && h_cnt <= 460 && v_cnt >= 100 && v_cnt <= 120) || (h_cnt >= 440 && h_cnt <= 460 && v_cnt >= 160 && v_cnt <= 180))
                                         {vgaRed, vgaGreen, vgaBlue} = 12'hfff; // bagel(in)
                                    else
                                        {vgaRed, vgaGreen, vgaBlue} = 12'hfde;
                                end
                                1'b1:begin
                                    if(!valid)
                                        {vgaRed, vgaGreen, vgaBlue} = 12'h0;
                                    else
                                        {vgaRed, vgaGreen, vgaBlue} = 12'hfde;
                                end
                            endcase    
			end
			3'b001:begin
				if(!valid)
					 {vgaRed, vgaGreen, vgaBlue} = 12'h0;
				else if(((h_cnt>=x+66&&h_cnt<x+72)&&(v_cnt>=370&&v_cnt<375))||((h_cnt>=x+54&&h_cnt<x+60)&&(v_cnt>=370&&v_cnt<380))||((h_cnt>=x+54&&h_cnt<x+78)&&(v_cnt>=390&&v_cnt<395))||((h_cnt>=x+60&&h_cnt<x+66)&&(v_cnt>=385&&v_cnt<390)))
					{vgaRed, vgaGreen, vgaBlue} = 12'h001;//BLACK
				else if(((h_cnt>=x+36&&h_cnt<x+42)&&(v_cnt>=400&&v_cnt<405))||((h_cnt>=x+60&&h_cnt<x+66)&&(v_cnt>=400&&v_cnt<405))||((h_cnt>=x+42&&h_cnt<x+48)&&(v_cnt>=405&&v_cnt<420))||((h_cnt>=x+48&&h_cnt<x+66)&&(v_cnt>=410&&v_cnt<415))||((h_cnt>=x+66&&h_cnt<x+72)&&(v_cnt>=405&&v_cnt<410))||((h_cnt>=x+72&&h_cnt<x+84)&&(v_cnt>=410&&v_cnt<425))||((h_cnt>=x+54&&h_cnt<x+72)&&(v_cnt>=415&&v_cnt<425))||((h_cnt>=x+24&&h_cnt<x+60)&&(v_cnt>=425&&v_cnt<430))||((h_cnt>=x+24&&h_cnt<x+54)&&(v_cnt>=420&&v_cnt<425))||((h_cnt>=x+24&&h_cnt<x+30)&&(v_cnt>=415&&v_cnt<420))||((h_cnt>=x+36&&h_cnt<x+42)&&(v_cnt>=415&&v_cnt<420)))
					{vgaRed, vgaGreen, vgaBlue} = 12'h00f;//BLUE
				else if(((h_cnt>=x+66&&h_cnt<x+72)&&(v_cnt>=410&&v_cnt<415))||((h_cnt>=x+48&&h_cnt<x+54)&&(v_cnt>=415&&v_cnt<420)))
					{vgaRed, vgaGreen, vgaBlue} = 12'hff0;//Y
				else if(((h_cnt>=x+90&&h_cnt<x+96)&&(v_cnt>=400&&v_cnt<425))||((h_cnt>=x+84&&h_cnt<x+90)&&(v_cnt>=405&&v_cnt<425))||((h_cnt>=x+18&&h_cnt<x+24)&&(v_cnt>=375&&v_cnt<405))||((h_cnt>=x+24&&h_cnt<x+42)&&(v_cnt>=370&&v_cnt<375))||((h_cnt>=x+30&&h_cnt<x+36)&&(v_cnt>=375&&v_cnt<390))||((h_cnt>=x+24&&h_cnt<x+30)&&(v_cnt>=390&&v_cnt<395))||((h_cnt>=x+36&&h_cnt<x+42)&&(v_cnt>=385&&v_cnt<390))||((h_cnt>=x+6&&h_cnt<x+18)&&(v_cnt>=425&&v_cnt<435))||((h_cnt>=x+12&&h_cnt<x+30)&&(v_cnt>=420&&v_cnt<425))||((h_cnt>=x+18&&h_cnt<x+24)&&(v_cnt>=425&&v_cnt<430)))
					{vgaRed, vgaGreen, vgaBlue} = 12'hfa2;              
				else if(((h_cnt>=x+72&&h_cnt<x+90)&&(v_cnt>=360&&v_cnt<365))||((h_cnt>=x+78&&h_cnt<x+90)&&(v_cnt>=365&&v_cnt<370))||((h_cnt>=x+60&&h_cnt<x+66)&&(v_cnt>=370&&v_cnt<395))||((h_cnt>=x+66&&h_cnt<x+72)&&(v_cnt>=375&&v_cnt<390))||((h_cnt>=x+72&&h_cnt<x+78)&&(v_cnt>=385&&v_cnt<390))||((h_cnt>=x+78&&h_cnt<x+84)&&(v_cnt>=385&&v_cnt<390))||((h_cnt>=x+30&&h_cnt<x+54)&&(v_cnt>=390&&v_cnt<400))||((h_cnt>=x+42&&h_cnt<x+54)&&(v_cnt>=370&&v_cnt<390))||((h_cnt>=x+24&&h_cnt<x+30)&&(v_cnt>=375&&v_cnt<390))||((h_cnt>=x+36&&h_cnt<x+42)&&(v_cnt>=375&&v_cnt<385))||((h_cnt>=x+54&&h_cnt<x+72)&&(v_cnt>=395&&v_cnt<400))||((h_cnt>=x+54&&h_cnt<x+60)&&(v_cnt>=380&&v_cnt<390))||((h_cnt>=x+0&&h_cnt<x+12)&&(v_cnt>=405&&v_cnt<415))||((h_cnt>=x+18&&h_cnt<x+24)&&(v_cnt>=410&&v_cnt<415))||((h_cnt>=x+6&&h_cnt<x+12)&&(v_cnt>=415&&v_cnt<420)))
					{vgaRed, vgaGreen, vgaBlue} = 12'hf70;
				else if(((h_cnt>=x+24&&h_cnt<x+78)&&(v_cnt>=365&&v_cnt<370))||((h_cnt>=x+30&&h_cnt<x+60)&&(v_cnt>=360&&v_cnt<365))||((h_cnt>=x+72&&h_cnt<x+90)&&(v_cnt>=370&&v_cnt<380))||((h_cnt>=x+12&&h_cnt<x+36)&&(v_cnt>=400&&v_cnt<410))||((h_cnt>=x+18&&h_cnt<x+42)&&(v_cnt>=405&&v_cnt<415))||((h_cnt>=x+42&&h_cnt<x+60)&&(v_cnt>=400&&v_cnt<405))||((h_cnt>=x+48&&h_cnt<x+66)&&(v_cnt>=405&&v_cnt<410))||((h_cnt>=x+78&&h_cnt<x+90)&&(v_cnt>=380&&v_cnt<385))||((h_cnt>=x+66&&h_cnt<x+78)&&(v_cnt>=400&&v_cnt<405))||((h_cnt>=x+72&&h_cnt<x+84)&&(v_cnt>=395&&v_cnt<400))||((h_cnt>=x+78&&h_cnt<x+84)&&(v_cnt>=390&&v_cnt<395))||((h_cnt>=x+30&&h_cnt<x+36)&&(v_cnt>=415&&v_cnt<420))||((h_cnt>=x+84&&h_cnt<x+90)&&(v_cnt>=385&&v_cnt<390)))
					{vgaRed, vgaGreen, vgaBlue} = 12'hf00;//red

				else if((h_cnt>=branch1_x+10 && h_cnt<branch1_x+12)&&(v_cnt>=branch1_y+8 && v_cnt<branch1_y+39) || (h_cnt>=branch1_x+7 && h_cnt<branch1_x+10 && v_cnt==branch1_y+10) || (h_cnt==branch1_x+6 && v_cnt>=branch1_y+8 && v_cnt<branch1_y+10) || (h_cnt==branch1_x+5 && v_cnt==branch1_y+8) || (h_cnt>=branch1_x+3 && h_cnt<branch1_x+5 && v_cnt==branch1_y+7) || (h_cnt==branch1_x+6 && v_cnt>=branch1_y+8 && v_cnt<branch1_y+10) || (h_cnt==branch1_x+2 && v_cnt>=branch1_y+5 && v_cnt<branch1_y+7) || (h_cnt==branch1_x+1 && v_cnt==branch1_y+5) || (h_cnt==branch1_x && v_cnt==branch1_y+4) || (h_cnt>=branch1_x+11 && h_cnt<branch1_x+14 && v_cnt==branch1_y+7) || (h_cnt>=branch1_x+14 && h_cnt<branch1_x+16 && v_cnt==branch1_y+5) || (h_cnt==branch1_x+14 && v_cnt==branch1_y+6) || (h_cnt>=branch1_x+16 && h_cnt<branch1_x+17 && v_cnt==branch1_y+4) || (h_cnt>=branch1_x+18 && h_cnt<branch1_x+19 && v_cnt==branch1_y+1) || (h_cnt==branch1_x+17 && v_cnt==branch1_y+3) || (h_cnt==branch1_x+18 && v_cnt==branch1_y+2))
					{vgaRed, vgaGreen, vgaBlue} = 12'h644; // brown
				else if((h_cnt>=branch1_x+5 && h_cnt<branch1_x+6 && v_cnt==branch1_y+10) || (h_cnt>=branch1_x+2 && h_cnt<branch1_x+4 && v_cnt==branch1_y+8) || (h_cnt>=branch1_x && h_cnt<branch1_x+1 && v_cnt==branch1_y+6) || (h_cnt>=branch1_x+3 && h_cnt<branch1_x+5 && v_cnt==branch1_y+6) || (h_cnt>=branch1_x+1 && h_cnt<branch1_x+2 && v_cnt==branch1_y+4) || (h_cnt>=branch1_x+13 && h_cnt<branch1_x+14 && v_cnt==branch1_y+4) || (h_cnt>=branch1_x+15 && h_cnt<branch1_x+16 && v_cnt==branch1_y+3) || (h_cnt>=branch1_x+16 && h_cnt<branch1_x+17 && v_cnt==branch1_y+5) || (h_cnt>=branch1_x+19 && h_cnt<branch1_x+20 && v_cnt==branch1_y) || (h_cnt==branch1_x+7 && v_cnt>=branch1_y+7 && v_cnt<branch1_y+8) || (h_cnt==branch1_x+17 && v_cnt>=branch1_y+1 && v_cnt<branch1_y+2) || (h_cnt==branch1_x+18 && v_cnt>=branch1_y+3 && v_cnt<branch1_y+4) || (h_cnt==branch1_x+2 && v_cnt==branch1_y+3) || (h_cnt==branch1_x+2 && v_cnt==branch1_y+7) || (h_cnt==branch1_x+4 && v_cnt==branch1_y+9) || (h_cnt==branch1_x+6 && v_cnt==branch1_y+11) || (h_cnt==branch1_x+12 && v_cnt==branch1_y+6) || (h_cnt==branch1_x+14 && v_cnt==branch1_y+8) || (h_cnt==branch1_x+19 && v_cnt==branch1_y+2) || (h_cnt==branch1_x+20 && v_cnt==branch1_y+1))
					{vgaRed, vgaGreen, vgaBlue} = 12'h9b2; // green

				else if((h_cnt>=branch2_x+10 && h_cnt<branch2_x+12)&&(v_cnt>=branch2_y+8 && v_cnt<branch2_y+39) || (h_cnt>=branch2_x+7 && h_cnt<branch2_x+10 && v_cnt==branch2_y+10) || (h_cnt==branch2_x+6 && v_cnt>=branch2_y+8 && v_cnt<branch2_y+10) || (h_cnt==branch2_x+5 && v_cnt==branch2_y+8) || (h_cnt>=branch2_x+3 && h_cnt<branch2_x+5 && v_cnt==branch2_y+7) || (h_cnt==branch2_x+6 && v_cnt>=branch2_y+8 && v_cnt<branch2_y+10) || (h_cnt==branch2_x+2 && v_cnt>=branch2_y+5 && v_cnt<branch2_y+7) || (h_cnt==branch2_x+1 && v_cnt==branch2_y+5) || (h_cnt==branch2_x && v_cnt==branch2_y+4) || (h_cnt>=branch2_x+11 && h_cnt<branch2_x+14 && v_cnt==branch2_y+7) || (h_cnt>=branch2_x+14 && h_cnt<branch2_x+16 && v_cnt==branch2_y+5) || (h_cnt==branch2_x+14 && v_cnt==branch2_y+6) || (h_cnt>=branch2_x+16 && h_cnt<branch2_x+17 && v_cnt==branch2_y+4) || (h_cnt>=branch2_x+18 && h_cnt<branch2_x+19 && v_cnt==branch2_y+1) || (h_cnt==branch2_x+17 && v_cnt==branch2_y+3) || (h_cnt==branch2_x+18 && v_cnt==branch2_y+2))
					{vgaRed, vgaGreen, vgaBlue} = 12'h644; // brown
				else if((h_cnt>=branch2_x+5 && h_cnt<branch2_x+6 && v_cnt==branch2_y+10) || (h_cnt>=branch2_x+2 && h_cnt<branch2_x+4 && v_cnt==branch2_y+8) || (h_cnt>=branch2_x && h_cnt<branch2_x+1 && v_cnt==branch2_y+6) || (h_cnt>=branch2_x+3 && h_cnt<branch2_x+5 && v_cnt==branch2_y+6) || (h_cnt>=branch2_x+1 && h_cnt<branch2_x+2 && v_cnt==branch2_y+4) || (h_cnt>=branch2_x+13 && h_cnt<branch2_x+14 && v_cnt==branch2_y+4) || (h_cnt>=branch2_x+15 && h_cnt<branch2_x+16 && v_cnt==branch2_y+3) || (h_cnt>=branch2_x+16 && h_cnt<branch2_x+17 && v_cnt==branch2_y+5) || (h_cnt>=branch2_x+19 && h_cnt<branch2_x+20 && v_cnt==branch2_y) || (h_cnt==branch2_x+7 && v_cnt>=branch2_y+7 && v_cnt<branch2_y+8) || (h_cnt==branch2_x+17 && v_cnt>=branch2_y+1 && v_cnt<branch2_y+2) || (h_cnt==branch2_x+18 && v_cnt>=branch2_y+3 && v_cnt<branch2_y+4) || (h_cnt==branch2_x+2 && v_cnt==branch2_y+3) || (h_cnt==branch2_x+2 && v_cnt==branch2_y+7) || (h_cnt==branch2_x+4 && v_cnt==branch2_y+9) || (h_cnt==branch2_x+6 && v_cnt==branch2_y+11) || (h_cnt==branch2_x+12 && v_cnt==branch2_y+6) || (h_cnt==branch2_x+14 && v_cnt==branch2_y+8) || (h_cnt==branch2_x+19 && v_cnt==branch2_y+2) || (h_cnt==branch2_x+20 && v_cnt==branch2_y+1))
					{vgaRed, vgaGreen, vgaBlue} = 12'h9b2; // green

				else if((h_cnt>=branch3_x+10 && h_cnt<branch3_x+12)&&(v_cnt>=branch3_y+8 && v_cnt<branch3_y+39) || (h_cnt>=branch3_x+7 && h_cnt<branch3_x+10 && v_cnt==branch3_y+10) || (h_cnt==branch3_x+6 && v_cnt>=branch3_y+8 && v_cnt<branch3_y+10) || (h_cnt==branch3_x+5 && v_cnt==branch3_y+8) || (h_cnt>=branch3_x+3 && h_cnt<branch3_x+5 && v_cnt==branch3_y+7) || (h_cnt==branch3_x+6 && v_cnt>=branch3_y+8 && v_cnt<branch3_y+10) || (h_cnt==branch3_x+2 && v_cnt>=branch3_y+5 && v_cnt<branch3_y+7) || (h_cnt==branch3_x+1 && v_cnt==branch3_y+5) || (h_cnt==branch3_x && v_cnt==branch3_y+4) || (h_cnt>=branch3_x+11 && h_cnt<branch3_x+14 && v_cnt==branch3_y+7) || (h_cnt>=branch3_x+14 && h_cnt<branch3_x+16 && v_cnt==branch3_y+5) || (h_cnt==branch3_x+14 && v_cnt==branch3_y+6) || (h_cnt>=branch3_x+16 && h_cnt<branch3_x+17 && v_cnt==branch3_y+4) || (h_cnt>=branch3_x+18 && h_cnt<branch3_x+19 && v_cnt==branch3_y+1) || (h_cnt==branch3_x+17 && v_cnt==branch3_y+3) || (h_cnt==branch3_x+18 && v_cnt==branch3_y+2))
					{vgaRed, vgaGreen, vgaBlue} = 12'h644; // brown
				else if((h_cnt>=branch3_x+5 && h_cnt<branch3_x+6 && v_cnt==branch3_y+10) || (h_cnt>=branch3_x+2 && h_cnt<branch3_x+4 && v_cnt==branch3_y+8) || (h_cnt>=branch3_x && h_cnt<branch3_x+1 && v_cnt==branch3_y+6) || (h_cnt>=branch3_x+3 && h_cnt<branch3_x+5 && v_cnt==branch3_y+6) || (h_cnt>=branch3_x+1 && h_cnt<branch3_x+2 && v_cnt==branch3_y+4) || (h_cnt>=branch3_x+13 && h_cnt<branch3_x+14 && v_cnt==branch3_y+4) || (h_cnt>=branch3_x+15 && h_cnt<branch3_x+16 && v_cnt==branch3_y+3) || (h_cnt>=branch3_x+16 && h_cnt<branch3_x+17 && v_cnt==branch3_y+5) || (h_cnt>=branch3_x+19 && h_cnt<branch3_x+20 && v_cnt==branch3_y) || (h_cnt==branch3_x+7 && v_cnt>=branch3_y+7 && v_cnt<branch3_y+8) || (h_cnt==branch3_x+17 && v_cnt>=branch3_y+1 && v_cnt<branch3_y+2) || (h_cnt==branch3_x+18 && v_cnt>=branch3_y+3 && v_cnt<branch3_y+4) || (h_cnt==branch3_x+2 && v_cnt==branch3_y+3) || (h_cnt==branch3_x+2 && v_cnt==branch3_y+7) || (h_cnt==branch3_x+4 && v_cnt==branch3_y+9) || (h_cnt==branch3_x+6 && v_cnt==branch3_y+11) || (h_cnt==branch3_x+12 && v_cnt==branch3_y+6) || (h_cnt==branch3_x+14 && v_cnt==branch3_y+8) || (h_cnt==branch3_x+19 && v_cnt==branch3_y+2) || (h_cnt==branch3_x+20 && v_cnt==branch3_y+1))
					{vgaRed, vgaGreen, vgaBlue} = 12'h9b2; // green

				else if((h_cnt>=branch4_x+10 && h_cnt<branch4_x+12)&&(v_cnt>=branch4_y+8 && v_cnt<branch4_y+39) || (h_cnt>=branch4_x+7 && h_cnt<branch4_x+10 && v_cnt==branch4_y+10) || (h_cnt==branch4_x+6 && v_cnt>=branch4_y+8 && v_cnt<branch4_y+10) || (h_cnt==branch4_x+5 && v_cnt==branch4_y+8) || (h_cnt>=branch4_x+3 && h_cnt<branch4_x+5 && v_cnt==branch4_y+7) || (h_cnt==branch4_x+6 && v_cnt>=branch4_y+8 && v_cnt<branch4_y+10) || (h_cnt==branch4_x+2 && v_cnt>=branch4_y+5 && v_cnt<branch4_y+7) || (h_cnt==branch4_x+1 && v_cnt==branch4_y+5) || (h_cnt==branch4_x && v_cnt==branch4_y+4) || (h_cnt>=branch4_x+11 && h_cnt<branch4_x+14 && v_cnt==branch4_y+7) || (h_cnt>=branch4_x+14 && h_cnt<branch4_x+16 && v_cnt==branch4_y+5) || (h_cnt==branch4_x+14 && v_cnt==branch4_y+6) || (h_cnt>=branch4_x+16 && h_cnt<branch4_x+17 && v_cnt==branch4_y+4) || (h_cnt>=branch4_x+18 && h_cnt<branch4_x+19 && v_cnt==branch4_y+1) || (h_cnt==branch4_x+17 && v_cnt==branch4_y+3) || (h_cnt==branch4_x+18 && v_cnt==branch4_y+2))
					{vgaRed, vgaGreen, vgaBlue} = 12'h644; // brown
				else if((h_cnt>=branch4_x+5 && h_cnt<branch4_x+6 && v_cnt==branch4_y+10) || (h_cnt>=branch4_x+2 && h_cnt<branch4_x+4 && v_cnt==branch4_y+8) || (h_cnt>=branch4_x && h_cnt<branch4_x+1 && v_cnt==branch4_y+6) || (h_cnt>=branch4_x+3 && h_cnt<branch4_x+5 && v_cnt==branch4_y+6) || (h_cnt>=branch4_x+1 && h_cnt<branch4_x+2 && v_cnt==branch4_y+4) || (h_cnt>=branch4_x+13 && h_cnt<branch4_x+14 && v_cnt==branch4_y+4) || (h_cnt>=branch4_x+15 && h_cnt<branch4_x+16 && v_cnt==branch4_y+3) || (h_cnt>=branch4_x+16 && h_cnt<branch4_x+17 && v_cnt==branch4_y+5) || (h_cnt>=branch4_x+19 && h_cnt<branch4_x+20 && v_cnt==branch4_y) || (h_cnt==branch4_x+7 && v_cnt>=branch4_y+7 && v_cnt<branch4_y+8) || (h_cnt==branch4_x+17 && v_cnt>=branch4_y+1 && v_cnt<branch4_y+2) || (h_cnt==branch4_x+18 && v_cnt>=branch4_y+3 && v_cnt<branch4_y+4) || (h_cnt==branch4_x+2 && v_cnt==branch4_y+3) || (h_cnt==branch4_x+2 && v_cnt==branch4_y+7) || (h_cnt==branch4_x+4 && v_cnt==branch4_y+9) || (h_cnt==branch4_x+6 && v_cnt==branch4_y+11) || (h_cnt==branch4_x+12 && v_cnt==branch4_y+6) || (h_cnt==branch4_x+14 && v_cnt==branch4_y+8) || (h_cnt==branch4_x+19 && v_cnt==branch4_y+2) || (h_cnt==branch4_x+20 && v_cnt==branch4_y+1))
					{vgaRed, vgaGreen, vgaBlue} = 12'h9b2; // green
					
				else if((h_cnt>=branch5_x+10 && h_cnt<branch5_x+12)&&(v_cnt>=branch5_y+8 && v_cnt<branch5_y+39) || (h_cnt>=branch5_x+7 && h_cnt<branch5_x+10 && v_cnt==branch5_y+10) || (h_cnt==branch5_x+6 && v_cnt>=branch5_y+8 && v_cnt<branch5_y+10) || (h_cnt==branch5_x+5 && v_cnt==branch5_y+8) || (h_cnt>=branch5_x+3 && h_cnt<branch5_x+5 && v_cnt==branch5_y+7) || (h_cnt==branch5_x+6 && v_cnt>=branch5_y+8 && v_cnt<branch5_y+10) || (h_cnt==branch5_x+2 && v_cnt>=branch5_y+5 && v_cnt<branch5_y+7) || (h_cnt==branch5_x+1 && v_cnt==branch5_y+5) || (h_cnt==branch5_x && v_cnt==branch5_y+4) || (h_cnt>=branch5_x+11 && h_cnt<branch5_x+14 && v_cnt==branch5_y+7) || (h_cnt>=branch5_x+14 && h_cnt<branch5_x+16 && v_cnt==branch5_y+5) || (h_cnt==branch5_x+14 && v_cnt==branch5_y+6) || (h_cnt>=branch5_x+16 && h_cnt<branch5_x+17 && v_cnt==branch5_y+4) || (h_cnt>=branch5_x+18 && h_cnt<branch5_x+19 && v_cnt==branch5_y+1) || (h_cnt==branch5_x+17 && v_cnt==branch5_y+3) || (h_cnt==branch5_x+18 && v_cnt==branch5_y+2))
					{vgaRed, vgaGreen, vgaBlue} = 12'h644; // brown
				else if((h_cnt>=branch5_x+5 && h_cnt<branch5_x+6 && v_cnt==branch5_y+10) || (h_cnt>=branch5_x+2 && h_cnt<branch5_x+4 && v_cnt==branch5_y+8) || (h_cnt>=branch5_x && h_cnt<branch5_x+1 && v_cnt==branch5_y+6) || (h_cnt>=branch5_x+3 && h_cnt<branch5_x+5 && v_cnt==branch5_y+6) || (h_cnt>=branch5_x+1 && h_cnt<branch5_x+2 && v_cnt==branch5_y+4) || (h_cnt>=branch5_x+13 && h_cnt<branch5_x+14 && v_cnt==branch5_y+4) || (h_cnt>=branch5_x+15 && h_cnt<branch5_x+16 && v_cnt==branch5_y+3) || (h_cnt>=branch5_x+16 && h_cnt<branch5_x+17 && v_cnt==branch5_y+5) || (h_cnt>=branch5_x+19 && h_cnt<branch5_x+20 && v_cnt==branch5_y) || (h_cnt==branch5_x+7 && v_cnt>=branch5_y+7 && v_cnt<branch5_y+8) || (h_cnt==branch5_x+17 && v_cnt>=branch5_y+1 && v_cnt<branch5_y+2) || (h_cnt==branch5_x+18 && v_cnt>=branch5_y+3 && v_cnt<branch5_y+4) || (h_cnt==branch5_x+2 && v_cnt==branch5_y+3) || (h_cnt==branch5_x+2 && v_cnt==branch5_y+7) || (h_cnt==branch5_x+4 && v_cnt==branch5_y+9) || (h_cnt==branch5_x+6 && v_cnt==branch5_y+11) || (h_cnt==branch5_x+12 && v_cnt==branch5_y+6) || (h_cnt==branch5_x+14 && v_cnt==branch5_y+8) || (h_cnt==branch5_x+19 && v_cnt==branch5_y+2) || (h_cnt==branch5_x+20 && v_cnt==branch5_y+1))
					{vgaRed, vgaGreen, vgaBlue} = 12'h9b2; // green
		
				else if((h_cnt >= bagel1_x+12 && h_cnt <= bagel1_x+26 && v_cnt >= bagel1_y && v_cnt <= bagel1_y+2)||(h_cnt >= bagel1_x+8 && h_cnt <= bagel1_x+12 && v_cnt >= bagel1_y+2 && v_cnt <= bagel1_y+4)||(h_cnt >= bagel1_x+26 && h_cnt <= bagel1_x+30 && v_cnt >= bagel1_y+2 && v_cnt <= bagel1_y+4)||(h_cnt >= bagel1_x+6 && h_cnt <= bagel1_x+8 && v_cnt >= bagel1_y+4 && v_cnt <= bagel1_y+6)||(h_cnt >= bagel1_x+30 && h_cnt <= bagel1_x+32 && v_cnt >= bagel1_y+4 && v_cnt <= bagel1_y+6)||(h_cnt >= bagel1_x+4 && h_cnt <= bagel1_x+6 && v_cnt >= bagel1_y+6 && v_cnt <= bagel1_y+8)||(h_cnt >= bagel1_x+32 && h_cnt <= bagel1_x+34 && v_cnt >= bagel1_y+6 && v_cnt <= bagel1_y+8)||(h_cnt >= bagel1_x+2 && h_cnt <= bagel1_x+4 && v_cnt >= bagel1_y+8 && v_cnt <= bagel1_y+12)||(h_cnt >= bagel1_x+34 && h_cnt <= bagel1_x+36 && v_cnt >= bagel1_y+8 && v_cnt <= bagel1_y+12)||(h_cnt >= bagel1_x && h_cnt <= bagel1_x+2 && v_cnt >= bagel1_y+12 && v_cnt <= bagel1_y+24)||(h_cnt >= bagel1_x+36 && h_cnt <= bagel1_x+38 && v_cnt >= bagel1_y+12 && v_cnt <= bagel1_y+24)||(h_cnt >= bagel1_x+2 && h_cnt <= bagel1_x+4 && v_cnt >= bagel1_y+24 && v_cnt <= bagel1_y+28)||(h_cnt >= bagel1_x+34 && h_cnt <= bagel1_x+36 && v_cnt >= bagel1_y+24 && v_cnt <= bagel1_y+28)||(h_cnt >= bagel1_x+4 && h_cnt <= bagel1_x+6 && v_cnt >= bagel1_y+28 && v_cnt <= bagel1_y+30)||(h_cnt >= bagel1_x+32 && h_cnt <= bagel1_x+34 && v_cnt >= bagel1_y+28 && v_cnt <= bagel1_y+30)||(h_cnt >= bagel1_x+6 && h_cnt <= bagel1_x+8 && v_cnt >= bagel1_y+30 && v_cnt <= bagel1_y+32)||(h_cnt >= bagel1_x+30 && h_cnt <= bagel1_x+32 && v_cnt >= bagel1_y+30 && v_cnt <= bagel1_y+32)||(h_cnt >= bagel1_x+8 && h_cnt <= bagel1_x+12 && v_cnt >= bagel1_y+32 && v_cnt <= bagel1_y+34)||(h_cnt >= bagel1_x+26 && h_cnt <= bagel1_x+30 && v_cnt >= bagel1_y+32 && v_cnt <= bagel1_y+34)||(h_cnt >= bagel1_x+12 && h_cnt <= bagel1_x+26 && v_cnt >= bagel1_y+34 && v_cnt <= bagel1_y+36)||(h_cnt >= bagel1_x+18 && h_cnt <= bagel1_x+22 && v_cnt >= bagel1_y+14 && v_cnt <= bagel1_y+16)||(h_cnt >= bagel1_x+18 && h_cnt <= bagel1_x+22 && v_cnt >= bagel1_y+20 && v_cnt <= bagel1_y+22)||(h_cnt >= bagel1_x+16 && h_cnt <= bagel1_x+18 && v_cnt >= bagel1_y+16 && v_cnt <= bagel1_y+20)||(h_cnt >= bagel1_x+22 && h_cnt <= bagel1_x+24 && v_cnt >= bagel1_y+16 && v_cnt <= bagel1_y+20))
					{vgaRed, vgaGreen, vgaBlue} = 12'h0; // black
				else if((h_cnt >= bagel1_x+14 && h_cnt <= bagel1_x+16 && v_cnt >= bagel1_y+2 && v_cnt <= bagel1_y+4)||(h_cnt >= bagel1_x+24 && h_cnt <= bagel1_x+26 && v_cnt >= bagel1_y+2 && v_cnt <= bagel1_y+4)||(h_cnt >= bagel1_x+8 && h_cnt <= bagel1_x+10 && v_cnt >= bagel1_y+4 && v_cnt <= bagel1_y+6)||(h_cnt >= bagel1_x+26 && h_cnt <= bagel1_x+28 && v_cnt >= bagel1_y+4 && v_cnt <= bagel1_y+6)||(h_cnt >= bagel1_x+6 && h_cnt <= bagel1_x+8 && v_cnt >= bagel1_y+6 && v_cnt <= bagel1_y+8)||(h_cnt >= bagel1_x+14 && h_cnt <= bagel1_x+26 && v_cnt >= bagel1_y+6 && v_cnt <= bagel1_y+8)||(h_cnt >= bagel1_x+28 && h_cnt <= bagel1_x+30 && v_cnt >= bagel1_y+6 && v_cnt <= bagel1_y+8)||(h_cnt >= bagel1_x+4 && h_cnt <= bagel1_x+6 && v_cnt >= bagel1_y+8 && v_cnt <= bagel1_y+10)||(h_cnt >= bagel1_x+12 && h_cnt <= bagel1_x+26 && v_cnt >= bagel1_y+8 && v_cnt <= bagel1_y+10)||(h_cnt >= bagel1_x+28 && h_cnt <= bagel1_x+32 && v_cnt >= bagel1_y+8 && v_cnt <= bagel1_y+10)||(h_cnt >= bagel1_x+10 && h_cnt <= bagel1_x+14 && v_cnt >= bagel1_y+10 && v_cnt <= bagel1_y+20)||(h_cnt >= bagel1_x+24 && h_cnt <= bagel1_x+26 && v_cnt >= bagel1_y+10 && v_cnt <= bagel1_y+14)||(h_cnt >= bagel1_x+30 && h_cnt <= bagel1_x+34 && v_cnt >= bagel1_y+10 && v_cnt <= bagel1_y+18)||(h_cnt >= bagel1_x+28 && h_cnt <= bagel1_x+32 && v_cnt >= bagel1_y+18 && v_cnt <= bagel1_y+20)||(h_cnt >= bagel1_x+4 && h_cnt <= bagel1_x+6 && v_cnt >= bagel1_y+18 && v_cnt <= bagel1_y+20)||(h_cnt >= bagel1_x+6 && h_cnt <= bagel1_x+10 && v_cnt >= bagel1_y+20 && v_cnt <= bagel1_y+22)||(h_cnt >= bagel1_x+12 && h_cnt <= bagel1_x+16 && v_cnt >= bagel1_y+20 && v_cnt <= bagel1_y+22)||(h_cnt >= bagel1_x+26 && h_cnt <= bagel1_x+30 && v_cnt >= bagel1_y+20 && v_cnt <= bagel1_y+22)||(h_cnt >= bagel1_x+34 && h_cnt <= bagel1_x+36 && v_cnt >= bagel1_y+20 && v_cnt <= bagel1_y+22)||(h_cnt >= bagel1_x+4 && h_cnt <= bagel1_x+6 && v_cnt >= bagel1_y+22 && v_cnt <= bagel1_y+24)||(h_cnt >= bagel1_x+8 && h_cnt <= bagel1_x+12 && v_cnt >= bagel1_y+22 && v_cnt <= bagel1_y+24)||(h_cnt >= bagel1_x+14 && h_cnt <= bagel1_x+22 && v_cnt >= bagel1_y+22 && v_cnt <= bagel1_y+24)||(h_cnt >= bagel1_x+24 && h_cnt <= bagel1_x+28 && v_cnt >= bagel1_y+22 && v_cnt <= bagel1_y+24)||(h_cnt >= bagel1_x+32 && h_cnt <= bagel1_x+34 && v_cnt >= bagel1_y+22 && v_cnt <= bagel1_y+24)||(h_cnt >= bagel1_x+6 && h_cnt <= bagel1_x+8 && v_cnt >= bagel1_y+24 && v_cnt <= bagel1_y+26)||(h_cnt >= bagel1_x+12 && h_cnt <= bagel1_x+24 && v_cnt >= bagel1_y+24 && v_cnt <= bagel1_y+26)||(h_cnt >= bagel1_x+30 && h_cnt <= bagel1_x+32 && v_cnt >= bagel1_y+24 && v_cnt <= bagel1_y+26)||(h_cnt >= bagel1_x+8 && h_cnt <= bagel1_x+10 && v_cnt >= bagel1_y+26 && v_cnt <= bagel1_y+28)||(h_cnt >= bagel1_x+28 && h_cnt <= bagel1_x+30 && v_cnt >= bagel1_y+26 && v_cnt <= bagel1_y+28)||(h_cnt >= bagel1_x+12 && h_cnt <= bagel1_x+14 && v_cnt >= bagel1_y+28 && v_cnt <= bagel1_y+30)||(h_cnt >= bagel1_x+24 && h_cnt <= bagel1_x+26 && v_cnt >= bagel1_y+28 && v_cnt <= bagel1_y+30))
					{vgaRed, vgaGreen, vgaBlue} = 12'hf9c; // baby pink
				else if((h_cnt >= bagel1_x+16 && h_cnt <= bagel1_x+24 && v_cnt >= bagel1_y+2 && v_cnt <= bagel1_y+4)||(h_cnt >= bagel1_x+10 && h_cnt <= bagel1_x+26 && v_cnt >= bagel1_y+4 && v_cnt <= bagel1_y+6)||(h_cnt >= bagel1_x+8 && h_cnt <= bagel1_x+14 && v_cnt >= bagel1_y+6 && v_cnt <= bagel1_y+8)||(h_cnt >= bagel1_x+26 && h_cnt <= bagel1_x+28 && v_cnt >= bagel1_y+6 && v_cnt <= bagel1_y+20)||(h_cnt >= bagel1_x+28 && h_cnt <= bagel1_x+30 && v_cnt >= bagel1_y+10 && v_cnt <= bagel1_y+18)||(h_cnt >= bagel1_x+24 && h_cnt <= bagel1_x+26 && v_cnt >= bagel1_y+14 && v_cnt <= bagel1_y+22)||(h_cnt >= bagel1_x+14 && h_cnt <= bagel1_x+24 && v_cnt >= bagel1_y+10 && v_cnt <= bagel1_y+14)||(h_cnt >= bagel1_x+4 && h_cnt <= bagel1_x+10 && v_cnt >= bagel1_y+10 && v_cnt <= bagel1_y+18)||(h_cnt >= bagel1_x+2 && h_cnt <= bagel1_x+4 && v_cnt >= bagel1_y+12 && v_cnt <= bagel1_y+24)||(h_cnt >= bagel1_x+6 && h_cnt <= bagel1_x+10 && v_cnt >= bagel1_y+18 && v_cnt <= bagel1_y+20)||(h_cnt >= bagel1_x+4 && h_cnt <= bagel1_x+6 && v_cnt >= bagel1_y+20 && v_cnt <= bagel1_y+22)||(h_cnt >= bagel1_x+34 && h_cnt <= bagel1_x+36 && v_cnt >= bagel1_y+12 && v_cnt <= bagel1_y+20)||(h_cnt >= bagel1_x+22 && h_cnt <= bagel1_x+24 && v_cnt >= bagel1_y+14 && v_cnt <= bagel1_y+16)||(h_cnt >= bagel1_x+14 && h_cnt <= bagel1_x+18 && v_cnt >= bagel1_y+14 && v_cnt <= bagel1_y+16)||(h_cnt >= bagel1_x+14 && h_cnt <= bagel1_x+16 && v_cnt >= bagel1_y+16 && v_cnt <= bagel1_y+20)||(h_cnt >= bagel1_x+32 && h_cnt <= bagel1_x+34 && v_cnt >= bagel1_y+18 && v_cnt <= bagel1_y+22)||(h_cnt >= bagel1_x+30 && h_cnt <= bagel1_x+32 && v_cnt >= bagel1_y+20 && v_cnt <= bagel1_y+24)||(h_cnt >= bagel1_x+28 && h_cnt <= bagel1_x+30 && v_cnt >= bagel1_y+22 && v_cnt <= bagel1_y+26)||(h_cnt >= bagel1_x+24 && h_cnt <= bagel1_x+28 && v_cnt >= bagel1_y+24 && v_cnt <= bagel1_y+28)||(h_cnt >= bagel1_x+14 && h_cnt <= bagel1_x+26 && v_cnt >= bagel1_y+26 && v_cnt <= bagel1_y+30)||(h_cnt >= bagel1_x+10 && h_cnt <= bagel1_x+14 && v_cnt >= bagel1_y+26 && v_cnt <= bagel1_y+28)||(h_cnt >= bagel1_x+8 && h_cnt <= bagel1_x+12 && v_cnt >= bagel1_y+24 && v_cnt <= bagel1_y+26)||(h_cnt >= bagel1_x+6 && h_cnt <= bagel1_x+12 && v_cnt >= bagel1_y+8 && v_cnt <= bagel1_y+10))
					{vgaRed, vgaGreen, vgaBlue} = 12'hf69; // light pink
				else if((h_cnt >= bagel1_x+12 && h_cnt <= bagel1_x+14 && v_cnt >= bagel1_y+2 && v_cnt <= bagel1_y+4)||(h_cnt >= bagel1_x+28 && h_cnt <= bagel1_x+30 && v_cnt >= bagel1_y+4 && v_cnt <= bagel1_y+6)||(h_cnt >= bagel1_x+30 && h_cnt <= bagel1_x+32 && v_cnt >= bagel1_y+6 && v_cnt <= bagel1_y+8)||(h_cnt >= bagel1_x+32 && h_cnt <= bagel1_x+34 && v_cnt >= bagel1_y+8 && v_cnt <= bagel1_y+10)||(h_cnt >= bagel1_x+10 && h_cnt <= bagel1_x+12 && v_cnt >= bagel1_y+20 && v_cnt <= bagel1_y+22)||(h_cnt >= bagel1_x+16 && h_cnt <= bagel1_x+18 && v_cnt >= bagel1_y+20 && v_cnt <= bagel1_y+22)||(h_cnt >= bagel1_x+22 && h_cnt <= bagel1_x+24 && v_cnt >= bagel1_y+20 && v_cnt <= bagel1_y+24)||(h_cnt >= bagel1_x+6 && h_cnt <= bagel1_x+8 && v_cnt >= bagel1_y+22 && v_cnt <= bagel1_y+24)||(h_cnt >= bagel1_x+32 && h_cnt <= bagel1_x+34 && v_cnt >= bagel1_y+24 && v_cnt <= bagel1_y+28)||(h_cnt >= bagel1_x+34 && h_cnt <= bagel1_x+36 && v_cnt >= bagel1_y+22 && v_cnt <= bagel1_y+24))
					{vgaRed, vgaGreen, vgaBlue} = 12'hf48; // dark pink
				else if((h_cnt >= bagel1_x+4 && h_cnt <= bagel1_x+6 && v_cnt >= bagel1_y+24 && v_cnt <= bagel1_y+28)||(h_cnt >= bagel1_x+6 && h_cnt <= bagel1_x+8 && v_cnt >= bagel1_y+26 && v_cnt <= bagel1_y+30)||(h_cnt >= bagel1_x+8 && h_cnt <= bagel1_x+12 && v_cnt >= bagel1_y+28 && v_cnt <= bagel1_y+32)||(h_cnt >= bagel1_x+12 && h_cnt <= bagel1_x+26 && v_cnt >= bagel1_y+30 && v_cnt <= bagel1_y+34)||(h_cnt >= bagel1_x+26 && h_cnt <= bagel1_x+30 && v_cnt >= bagel1_y+28 && v_cnt <= bagel1_y+32)||(h_cnt >= bagel1_x+30 && h_cnt <= bagel1_x+32 && v_cnt >= bagel1_y+26 && v_cnt <= bagel1_y+30)||(h_cnt >= bagel1_x+4 && h_cnt <= bagel1_x+6 && v_cnt >= bagel1_y+24 && v_cnt <= bagel1_y+28)||(h_cnt >= bagel1_x+12 && h_cnt <= bagel1_x+14 && v_cnt >= bagel1_y+22 && v_cnt <= bagel1_y+24))
					{vgaRed, vgaGreen, vgaBlue} = 12'hfd5; // yellow
				
				else if((h_cnt >= bagel2_x+12 && h_cnt <= bagel2_x+26 && v_cnt >= bagel2_y && v_cnt <= bagel2_y+2)||(h_cnt >= bagel2_x+8 && h_cnt <= bagel2_x+12 && v_cnt >= bagel2_y+2 && v_cnt <= bagel2_y+4)||(h_cnt >= bagel2_x+26 && h_cnt <= bagel2_x+30 && v_cnt >= bagel2_y+2 && v_cnt <= bagel2_y+4)||(h_cnt >= bagel2_x+6 && h_cnt <= bagel2_x+8 && v_cnt >= bagel2_y+4 && v_cnt <= bagel2_y+6)||(h_cnt >= bagel2_x+30 && h_cnt <= bagel2_x+32 && v_cnt >= bagel2_y+4 && v_cnt <= bagel2_y+6)||(h_cnt >= bagel2_x+4 && h_cnt <= bagel2_x+6 && v_cnt >= bagel2_y+6 && v_cnt <= bagel2_y+8)||(h_cnt >= bagel2_x+32 && h_cnt <= bagel2_x+34 && v_cnt >= bagel2_y+6 && v_cnt <= bagel2_y+8)||(h_cnt >= bagel2_x+2 && h_cnt <= bagel2_x+4 && v_cnt >= bagel2_y+8 && v_cnt <= bagel2_y+12)||(h_cnt >= bagel2_x+34 && h_cnt <= bagel2_x+36 && v_cnt >= bagel2_y+8 && v_cnt <= bagel2_y+12)||(h_cnt >= bagel2_x && h_cnt <= bagel2_x+2 && v_cnt >= bagel2_y+12 && v_cnt <= bagel2_y+24)||(h_cnt >= bagel2_x+36 && h_cnt <= bagel2_x+38 && v_cnt >= bagel2_y+12 && v_cnt <= bagel2_y+24)||(h_cnt >= bagel2_x+2 && h_cnt <= bagel2_x+4 && v_cnt >= bagel2_y+24 && v_cnt <= bagel2_y+28)||(h_cnt >= bagel2_x+34 && h_cnt <= bagel2_x+36 && v_cnt >= bagel2_y+24 && v_cnt <= bagel2_y+28)||(h_cnt >= bagel2_x+4 && h_cnt <= bagel2_x+6 && v_cnt >= bagel2_y+28 && v_cnt <= bagel2_y+30)||(h_cnt >= bagel2_x+32 && h_cnt <= bagel2_x+34 && v_cnt >= bagel2_y+28 && v_cnt <= bagel2_y+30)||(h_cnt >= bagel2_x+6 && h_cnt <= bagel2_x+8 && v_cnt >= bagel2_y+30 && v_cnt <= bagel2_y+32)||(h_cnt >= bagel2_x+30 && h_cnt <= bagel2_x+32 && v_cnt >= bagel2_y+30 && v_cnt <= bagel2_y+32)||(h_cnt >= bagel2_x+8 && h_cnt <= bagel2_x+12 && v_cnt >= bagel2_y+32 && v_cnt <= bagel2_y+34)||(h_cnt >= bagel2_x+26 && h_cnt <= bagel2_x+30 && v_cnt >= bagel2_y+32 && v_cnt <= bagel2_y+34)||(h_cnt >= bagel2_x+12 && h_cnt <= bagel2_x+26 && v_cnt >= bagel2_y+34 && v_cnt <= bagel2_y+36)||(h_cnt >= bagel2_x+18 && h_cnt <= bagel2_x+22 && v_cnt >= bagel2_y+14 && v_cnt <= bagel2_y+16)||(h_cnt >= bagel2_x+18 && h_cnt <= bagel2_x+22 && v_cnt >= bagel2_y+20 && v_cnt <= bagel2_y+22)||(h_cnt >= bagel2_x+16 && h_cnt <= bagel2_x+18 && v_cnt >= bagel2_y+16 && v_cnt <= bagel2_y+20)||(h_cnt >= bagel2_x+22 && h_cnt <= bagel2_x+24 && v_cnt >= bagel2_y+16 && v_cnt <= bagel2_y+20))
					{vgaRed, vgaGreen, vgaBlue} = 12'h0; // black
				else if((h_cnt >= bagel2_x+14 && h_cnt <= bagel2_x+16 && v_cnt >= bagel2_y+2 && v_cnt <= bagel2_y+4)||(h_cnt >= bagel2_x+24 && h_cnt <= bagel2_x+26 && v_cnt >= bagel2_y+2 && v_cnt <= bagel2_y+4)||(h_cnt >= bagel2_x+8 && h_cnt <= bagel2_x+10 && v_cnt >= bagel2_y+4 && v_cnt <= bagel2_y+6)||(h_cnt >= bagel2_x+26 && h_cnt <= bagel2_x+28 && v_cnt >= bagel2_y+4 && v_cnt <= bagel2_y+6)||(h_cnt >= bagel2_x+6 && h_cnt <= bagel2_x+8 && v_cnt >= bagel2_y+6 && v_cnt <= bagel2_y+8)||(h_cnt >= bagel2_x+14 && h_cnt <= bagel2_x+26 && v_cnt >= bagel2_y+6 && v_cnt <= bagel2_y+8)||(h_cnt >= bagel2_x+28 && h_cnt <= bagel2_x+30 && v_cnt >= bagel2_y+6 && v_cnt <= bagel2_y+8)||(h_cnt >= bagel2_x+4 && h_cnt <= bagel2_x+6 && v_cnt >= bagel2_y+8 && v_cnt <= bagel2_y+10)||(h_cnt >= bagel2_x+12 && h_cnt <= bagel2_x+26 && v_cnt >= bagel2_y+8 && v_cnt <= bagel2_y+10)||(h_cnt >= bagel2_x+28 && h_cnt <= bagel2_x+32 && v_cnt >= bagel2_y+8 && v_cnt <= bagel2_y+10)||(h_cnt >= bagel2_x+10 && h_cnt <= bagel2_x+14 && v_cnt >= bagel2_y+10 && v_cnt <= bagel2_y+20)||(h_cnt >= bagel2_x+24 && h_cnt <= bagel2_x+26 && v_cnt >= bagel2_y+10 && v_cnt <= bagel2_y+14)||(h_cnt >= bagel2_x+30 && h_cnt <= bagel2_x+34 && v_cnt >= bagel2_y+10 && v_cnt <= bagel2_y+18)||(h_cnt >= bagel2_x+28 && h_cnt <= bagel2_x+32 && v_cnt >= bagel2_y+18 && v_cnt <= bagel2_y+20)||(h_cnt >= bagel2_x+4 && h_cnt <= bagel2_x+6 && v_cnt >= bagel2_y+18 && v_cnt <= bagel2_y+20)||(h_cnt >= bagel2_x+6 && h_cnt <= bagel2_x+10 && v_cnt >= bagel2_y+20 && v_cnt <= bagel2_y+22)||(h_cnt >= bagel2_x+12 && h_cnt <= bagel2_x+16 && v_cnt >= bagel2_y+20 && v_cnt <= bagel2_y+22)||(h_cnt >= bagel2_x+26 && h_cnt <= bagel2_x+30 && v_cnt >= bagel2_y+20 && v_cnt <= bagel2_y+22)||(h_cnt >= bagel2_x+34 && h_cnt <= bagel2_x+36 && v_cnt >= bagel2_y+20 && v_cnt <= bagel2_y+22)||(h_cnt >= bagel2_x+4 && h_cnt <= bagel2_x+6 && v_cnt >= bagel2_y+22 && v_cnt <= bagel2_y+24)||(h_cnt >= bagel2_x+8 && h_cnt <= bagel2_x+12 && v_cnt >= bagel2_y+22 && v_cnt <= bagel2_y+24)||(h_cnt >= bagel2_x+14 && h_cnt <= bagel2_x+22 && v_cnt >= bagel2_y+22 && v_cnt <= bagel2_y+24)||(h_cnt >= bagel2_x+24 && h_cnt <= bagel2_x+28 && v_cnt >= bagel2_y+22 && v_cnt <= bagel2_y+24)||(h_cnt >= bagel2_x+32 && h_cnt <= bagel2_x+34 && v_cnt >= bagel2_y+22 && v_cnt <= bagel2_y+24)||(h_cnt >= bagel2_x+6 && h_cnt <= bagel2_x+8 && v_cnt >= bagel2_y+24 && v_cnt <= bagel2_y+26)||(h_cnt >= bagel2_x+12 && h_cnt <= bagel2_x+24 && v_cnt >= bagel2_y+24 && v_cnt <= bagel2_y+26)||(h_cnt >= bagel2_x+30 && h_cnt <= bagel2_x+32 && v_cnt >= bagel2_y+24 && v_cnt <= bagel2_y+26)||(h_cnt >= bagel2_x+8 && h_cnt <= bagel2_x+10 && v_cnt >= bagel2_y+26 && v_cnt <= bagel2_y+28)||(h_cnt >= bagel2_x+28 && h_cnt <= bagel2_x+30 && v_cnt >= bagel2_y+26 && v_cnt <= bagel2_y+28)||(h_cnt >= bagel2_x+12 && h_cnt <= bagel2_x+14 && v_cnt >= bagel2_y+28 && v_cnt <= bagel2_y+30)||(h_cnt >= bagel2_x+24 && h_cnt <= bagel2_x+26 && v_cnt >= bagel2_y+28 && v_cnt <= bagel2_y+30))
					{vgaRed, vgaGreen, vgaBlue} = 12'hf9c; // baby pink
				else if((h_cnt >= bagel2_x+16 && h_cnt <= bagel2_x+24 && v_cnt >= bagel2_y+2 && v_cnt <= bagel2_y+4)||(h_cnt >= bagel2_x+10 && h_cnt <= bagel2_x+26 && v_cnt >= bagel2_y+4 && v_cnt <= bagel2_y+6)||(h_cnt >= bagel2_x+8 && h_cnt <= bagel2_x+14 && v_cnt >= bagel2_y+6 && v_cnt <= bagel2_y+8)||(h_cnt >= bagel2_x+26 && h_cnt <= bagel2_x+28 && v_cnt >= bagel2_y+6 && v_cnt <= bagel2_y+20)||(h_cnt >= bagel2_x+28 && h_cnt <= bagel2_x+30 && v_cnt >= bagel2_y+10 && v_cnt <= bagel2_y+18)||(h_cnt >= bagel2_x+24 && h_cnt <= bagel2_x+26 && v_cnt >= bagel2_y+14 && v_cnt <= bagel2_y+22)||(h_cnt >= bagel2_x+14 && h_cnt <= bagel2_x+24 && v_cnt >= bagel2_y+10 && v_cnt <= bagel2_y+14)||(h_cnt >= bagel2_x+4 && h_cnt <= bagel2_x+10 && v_cnt >= bagel2_y+10 && v_cnt <= bagel2_y+18)||(h_cnt >= bagel2_x+2 && h_cnt <= bagel2_x+4 && v_cnt >= bagel2_y+12 && v_cnt <= bagel2_y+24)||(h_cnt >= bagel2_x+6 && h_cnt <= bagel2_x+10 && v_cnt >= bagel2_y+18 && v_cnt <= bagel2_y+20)||(h_cnt >= bagel2_x+4 && h_cnt <= bagel2_x+6 && v_cnt >= bagel2_y+20 && v_cnt <= bagel2_y+22)||(h_cnt >= bagel2_x+34 && h_cnt <= bagel2_x+36 && v_cnt >= bagel2_y+12 && v_cnt <= bagel2_y+20)||(h_cnt >= bagel2_x+22 && h_cnt <= bagel2_x+24 && v_cnt >= bagel2_y+14 && v_cnt <= bagel2_y+16)||(h_cnt >= bagel2_x+14 && h_cnt <= bagel2_x+18 && v_cnt >= bagel2_y+14 && v_cnt <= bagel2_y+16)||(h_cnt >= bagel2_x+14 && h_cnt <= bagel2_x+16 && v_cnt >= bagel2_y+16 && v_cnt <= bagel2_y+20)||(h_cnt >= bagel2_x+32 && h_cnt <= bagel2_x+34 && v_cnt >= bagel2_y+18 && v_cnt <= bagel2_y+22)||(h_cnt >= bagel2_x+30 && h_cnt <= bagel2_x+32 && v_cnt >= bagel2_y+20 && v_cnt <= bagel2_y+24)||(h_cnt >= bagel2_x+28 && h_cnt <= bagel2_x+30 && v_cnt >= bagel2_y+22 && v_cnt <= bagel2_y+26)||(h_cnt >= bagel2_x+24 && h_cnt <= bagel2_x+28 && v_cnt >= bagel2_y+24 && v_cnt <= bagel2_y+28)||(h_cnt >= bagel2_x+14 && h_cnt <= bagel2_x+26 && v_cnt >= bagel2_y+26 && v_cnt <= bagel2_y+30)||(h_cnt >= bagel2_x+10 && h_cnt <= bagel2_x+14 && v_cnt >= bagel2_y+26 && v_cnt <= bagel2_y+28)||(h_cnt >= bagel2_x+8 && h_cnt <= bagel2_x+12 && v_cnt >= bagel2_y+24 && v_cnt <= bagel2_y+26)||(h_cnt >= bagel2_x+6 && h_cnt <= bagel2_x+12 && v_cnt >= bagel2_y+8 && v_cnt <= bagel2_y+10))
					{vgaRed, vgaGreen, vgaBlue} = 12'hf69; // light pink
				else if((h_cnt >= bagel2_x+12 && h_cnt <= bagel2_x+14 && v_cnt >= bagel2_y+2 && v_cnt <= bagel2_y+4)||(h_cnt >= bagel2_x+28 && h_cnt <= bagel2_x+30 && v_cnt >= bagel2_y+4 && v_cnt <= bagel2_y+6)||(h_cnt >= bagel2_x+30 && h_cnt <= bagel2_x+32 && v_cnt >= bagel2_y+6 && v_cnt <= bagel2_y+8)||(h_cnt >= bagel2_x+32 && h_cnt <= bagel2_x+34 && v_cnt >= bagel2_y+8 && v_cnt <= bagel2_y+10)||(h_cnt >= bagel2_x+10 && h_cnt <= bagel2_x+12 && v_cnt >= bagel2_y+20 && v_cnt <= bagel2_y+22)||(h_cnt >= bagel2_x+16 && h_cnt <= bagel2_x+18 && v_cnt >= bagel2_y+20 && v_cnt <= bagel2_y+22)||(h_cnt >= bagel2_x+22 && h_cnt <= bagel2_x+24 && v_cnt >= bagel2_y+20 && v_cnt <= bagel2_y+24)||(h_cnt >= bagel2_x+6 && h_cnt <= bagel2_x+8 && v_cnt >= bagel2_y+22 && v_cnt <= bagel2_y+24)||(h_cnt >= bagel2_x+32 && h_cnt <= bagel2_x+34 && v_cnt >= bagel2_y+24 && v_cnt <= bagel2_y+28)||(h_cnt >= bagel2_x+34 && h_cnt <= bagel2_x+36 && v_cnt >= bagel2_y+22 && v_cnt <= bagel2_y+24))
					{vgaRed, vgaGreen, vgaBlue} = 12'hf48; // dark pink
				else if((h_cnt >= bagel2_x+4 && h_cnt <= bagel2_x+6 && v_cnt >= bagel2_y+24 && v_cnt <= bagel2_y+28)||(h_cnt >= bagel2_x+6 && h_cnt <= bagel2_x+8 && v_cnt >= bagel2_y+26 && v_cnt <= bagel2_y+30)||(h_cnt >= bagel2_x+8 && h_cnt <= bagel2_x+12 && v_cnt >= bagel2_y+28 && v_cnt <= bagel2_y+32)||(h_cnt >= bagel2_x+12 && h_cnt <= bagel2_x+26 && v_cnt >= bagel2_y+30 && v_cnt <= bagel2_y+34)||(h_cnt >= bagel2_x+26 && h_cnt <= bagel2_x+30 && v_cnt >= bagel2_y+28 && v_cnt <= bagel2_y+32)||(h_cnt >= bagel2_x+30 && h_cnt <= bagel2_x+32 && v_cnt >= bagel2_y+26 && v_cnt <= bagel2_y+30)||(h_cnt >= bagel2_x+4 && h_cnt <= bagel2_x+6 && v_cnt >= bagel2_y+24 && v_cnt <= bagel2_y+28)||(h_cnt >= bagel2_x+12 && h_cnt <= bagel2_x+14 && v_cnt >= bagel2_y+22 && v_cnt <= bagel2_y+24))
					{vgaRed, vgaGreen, vgaBlue} = 12'hfd5; // yellow
				
				else if((h_cnt >= bagel3_x+12 && h_cnt <= bagel3_x+26 && v_cnt >= bagel3_y && v_cnt <= bagel3_y+2)||(h_cnt >= bagel3_x+8 && h_cnt <= bagel3_x+12 && v_cnt >= bagel3_y+2 && v_cnt <= bagel3_y+4)||(h_cnt >= bagel3_x+26 && h_cnt <= bagel3_x+30 && v_cnt >= bagel3_y+2 && v_cnt <= bagel3_y+4)||(h_cnt >= bagel3_x+6 && h_cnt <= bagel3_x+8 && v_cnt >= bagel3_y+4 && v_cnt <= bagel3_y+6)||(h_cnt >= bagel3_x+30 && h_cnt <= bagel3_x+32 && v_cnt >= bagel3_y+4 && v_cnt <= bagel3_y+6)||(h_cnt >= bagel3_x+4 && h_cnt <= bagel3_x+6 && v_cnt >= bagel3_y+6 && v_cnt <= bagel3_y+8)||(h_cnt >= bagel3_x+32 && h_cnt <= bagel3_x+34 && v_cnt >= bagel3_y+6 && v_cnt <= bagel3_y+8)||(h_cnt >= bagel3_x+2 && h_cnt <= bagel3_x+4 && v_cnt >= bagel3_y+8 && v_cnt <= bagel3_y+12)||(h_cnt >= bagel3_x+34 && h_cnt <= bagel3_x+36 && v_cnt >= bagel3_y+8 && v_cnt <= bagel3_y+12)||(h_cnt >= bagel3_x && h_cnt <= bagel3_x+2 && v_cnt >= bagel3_y+12 && v_cnt <= bagel3_y+24)||(h_cnt >= bagel3_x+36 && h_cnt <= bagel3_x+38 && v_cnt >= bagel3_y+12 && v_cnt <= bagel3_y+24)||(h_cnt >= bagel3_x+2 && h_cnt <= bagel3_x+4 && v_cnt >= bagel3_y+24 && v_cnt <= bagel3_y+28)||(h_cnt >= bagel3_x+34 && h_cnt <= bagel3_x+36 && v_cnt >= bagel3_y+24 && v_cnt <= bagel3_y+28)||(h_cnt >= bagel3_x+4 && h_cnt <= bagel3_x+6 && v_cnt >= bagel3_y+28 && v_cnt <= bagel3_y+30)||(h_cnt >= bagel3_x+32 && h_cnt <= bagel3_x+34 && v_cnt >= bagel3_y+28 && v_cnt <= bagel3_y+30)||(h_cnt >= bagel3_x+6 && h_cnt <= bagel3_x+8 && v_cnt >= bagel3_y+30 && v_cnt <= bagel3_y+32)||(h_cnt >= bagel3_x+30 && h_cnt <= bagel3_x+32 && v_cnt >= bagel3_y+30 && v_cnt <= bagel3_y+32)||(h_cnt >= bagel3_x+8 && h_cnt <= bagel3_x+12 && v_cnt >= bagel3_y+32 && v_cnt <= bagel3_y+34)||(h_cnt >= bagel3_x+26 && h_cnt <= bagel3_x+30 && v_cnt >= bagel3_y+32 && v_cnt <= bagel3_y+34)||(h_cnt >= bagel3_x+12 && h_cnt <= bagel3_x+26 && v_cnt >= bagel3_y+34 && v_cnt <= bagel3_y+36)||(h_cnt >= bagel3_x+18 && h_cnt <= bagel3_x+22 && v_cnt >= bagel3_y+14 && v_cnt <= bagel3_y+16)||(h_cnt >= bagel3_x+18 && h_cnt <= bagel3_x+22 && v_cnt >= bagel3_y+20 && v_cnt <= bagel3_y+22)||(h_cnt >= bagel3_x+16 && h_cnt <= bagel3_x+18 && v_cnt >= bagel3_y+16 && v_cnt <= bagel3_y+20)||(h_cnt >= bagel3_x+22 && h_cnt <= bagel3_x+24 && v_cnt >= bagel3_y+16 && v_cnt <= bagel3_y+20))
					{vgaRed, vgaGreen, vgaBlue} = 12'h0; // black
				else if((h_cnt >= bagel3_x+14 && h_cnt <= bagel3_x+16 && v_cnt >= bagel3_y+2 && v_cnt <= bagel3_y+4)||(h_cnt >= bagel3_x+24 && h_cnt <= bagel3_x+26 && v_cnt >= bagel3_y+2 && v_cnt <= bagel3_y+4)||(h_cnt >= bagel3_x+8 && h_cnt <= bagel3_x+10 && v_cnt >= bagel3_y+4 && v_cnt <= bagel3_y+6)||(h_cnt >= bagel3_x+26 && h_cnt <= bagel3_x+28 && v_cnt >= bagel3_y+4 && v_cnt <= bagel3_y+6)||(h_cnt >= bagel3_x+6 && h_cnt <= bagel3_x+8 && v_cnt >= bagel3_y+6 && v_cnt <= bagel3_y+8)||(h_cnt >= bagel3_x+14 && h_cnt <= bagel3_x+26 && v_cnt >= bagel3_y+6 && v_cnt <= bagel3_y+8)||(h_cnt >= bagel3_x+28 && h_cnt <= bagel3_x+30 && v_cnt >= bagel3_y+6 && v_cnt <= bagel3_y+8)||(h_cnt >= bagel3_x+4 && h_cnt <= bagel3_x+6 && v_cnt >= bagel3_y+8 && v_cnt <= bagel3_y+10)||(h_cnt >= bagel3_x+12 && h_cnt <= bagel3_x+26 && v_cnt >= bagel3_y+8 && v_cnt <= bagel3_y+10)||(h_cnt >= bagel3_x+28 && h_cnt <= bagel3_x+32 && v_cnt >= bagel3_y+8 && v_cnt <= bagel3_y+10)||(h_cnt >= bagel3_x+10 && h_cnt <= bagel3_x+14 && v_cnt >= bagel3_y+10 && v_cnt <= bagel3_y+20)||(h_cnt >= bagel3_x+24 && h_cnt <= bagel3_x+26 && v_cnt >= bagel3_y+10 && v_cnt <= bagel3_y+14)||(h_cnt >= bagel3_x+30 && h_cnt <= bagel3_x+34 && v_cnt >= bagel3_y+10 && v_cnt <= bagel3_y+18)||(h_cnt >= bagel3_x+28 && h_cnt <= bagel3_x+32 && v_cnt >= bagel3_y+18 && v_cnt <= bagel3_y+20)||(h_cnt >= bagel3_x+4 && h_cnt <= bagel3_x+6 && v_cnt >= bagel3_y+18 && v_cnt <= bagel3_y+20)||(h_cnt >= bagel3_x+6 && h_cnt <= bagel3_x+10 && v_cnt >= bagel3_y+20 && v_cnt <= bagel3_y+22)||(h_cnt >= bagel3_x+12 && h_cnt <= bagel3_x+16 && v_cnt >= bagel3_y+20 && v_cnt <= bagel3_y+22)||(h_cnt >= bagel3_x+26 && h_cnt <= bagel3_x+30 && v_cnt >= bagel3_y+20 && v_cnt <= bagel3_y+22)||(h_cnt >= bagel3_x+34 && h_cnt <= bagel3_x+36 && v_cnt >= bagel3_y+20 && v_cnt <= bagel3_y+22)||(h_cnt >= bagel3_x+4 && h_cnt <= bagel3_x+6 && v_cnt >= bagel3_y+22 && v_cnt <= bagel3_y+24)||(h_cnt >= bagel3_x+8 && h_cnt <= bagel3_x+12 && v_cnt >= bagel3_y+22 && v_cnt <= bagel3_y+24)||(h_cnt >= bagel3_x+14 && h_cnt <= bagel3_x+22 && v_cnt >= bagel3_y+22 && v_cnt <= bagel3_y+24)||(h_cnt >= bagel3_x+24 && h_cnt <= bagel3_x+28 && v_cnt >= bagel3_y+22 && v_cnt <= bagel3_y+24)||(h_cnt >= bagel3_x+32 && h_cnt <= bagel3_x+34 && v_cnt >= bagel3_y+22 && v_cnt <= bagel3_y+24)||(h_cnt >= bagel3_x+6 && h_cnt <= bagel3_x+8 && v_cnt >= bagel3_y+24 && v_cnt <= bagel3_y+26)||(h_cnt >= bagel3_x+12 && h_cnt <= bagel3_x+24 && v_cnt >= bagel3_y+24 && v_cnt <= bagel3_y+26)||(h_cnt >= bagel3_x+30 && h_cnt <= bagel3_x+32 && v_cnt >= bagel3_y+24 && v_cnt <= bagel3_y+26)||(h_cnt >= bagel3_x+8 && h_cnt <= bagel3_x+10 && v_cnt >= bagel3_y+26 && v_cnt <= bagel3_y+28)||(h_cnt >= bagel3_x+28 && h_cnt <= bagel3_x+30 && v_cnt >= bagel3_y+26 && v_cnt <= bagel3_y+28)||(h_cnt >= bagel3_x+12 && h_cnt <= bagel3_x+14 && v_cnt >= bagel3_y+28 && v_cnt <= bagel3_y+30)||(h_cnt >= bagel3_x+24 && h_cnt <= bagel3_x+26 && v_cnt >= bagel3_y+28 && v_cnt <= bagel3_y+30))
					{vgaRed, vgaGreen, vgaBlue} = 12'hf9c; // baby pink
				else if((h_cnt >= bagel3_x+16 && h_cnt <= bagel3_x+24 && v_cnt >= bagel3_y+2 && v_cnt <= bagel3_y+4)||(h_cnt >= bagel3_x+10 && h_cnt <= bagel3_x+26 && v_cnt >= bagel3_y+4 && v_cnt <= bagel3_y+6)||(h_cnt >= bagel3_x+8 && h_cnt <= bagel3_x+14 && v_cnt >= bagel3_y+6 && v_cnt <= bagel3_y+8)||(h_cnt >= bagel3_x+26 && h_cnt <= bagel3_x+28 && v_cnt >= bagel3_y+6 && v_cnt <= bagel3_y+20)||(h_cnt >= bagel3_x+28 && h_cnt <= bagel3_x+30 && v_cnt >= bagel3_y+10 && v_cnt <= bagel3_y+18)||(h_cnt >= bagel3_x+24 && h_cnt <= bagel3_x+26 && v_cnt >= bagel3_y+14 && v_cnt <= bagel3_y+22)||(h_cnt >= bagel3_x+14 && h_cnt <= bagel3_x+24 && v_cnt >= bagel3_y+10 && v_cnt <= bagel3_y+14)||(h_cnt >= bagel3_x+4 && h_cnt <= bagel3_x+10 && v_cnt >= bagel3_y+10 && v_cnt <= bagel3_y+18)||(h_cnt >= bagel3_x+2 && h_cnt <= bagel3_x+4 && v_cnt >= bagel3_y+12 && v_cnt <= bagel3_y+24)||(h_cnt >= bagel3_x+6 && h_cnt <= bagel3_x+10 && v_cnt >= bagel3_y+18 && v_cnt <= bagel3_y+20)||(h_cnt >= bagel3_x+4 && h_cnt <= bagel3_x+6 && v_cnt >= bagel3_y+20 && v_cnt <= bagel3_y+22)||(h_cnt >= bagel3_x+34 && h_cnt <= bagel3_x+36 && v_cnt >= bagel3_y+12 && v_cnt <= bagel3_y+20)||(h_cnt >= bagel3_x+22 && h_cnt <= bagel3_x+24 && v_cnt >= bagel3_y+14 && v_cnt <= bagel3_y+16)||(h_cnt >= bagel3_x+14 && h_cnt <= bagel3_x+18 && v_cnt >= bagel3_y+14 && v_cnt <= bagel3_y+16)||(h_cnt >= bagel3_x+14 && h_cnt <= bagel3_x+16 && v_cnt >= bagel3_y+16 && v_cnt <= bagel3_y+20)||(h_cnt >= bagel3_x+32 && h_cnt <= bagel3_x+34 && v_cnt >= bagel3_y+18 && v_cnt <= bagel3_y+22)||(h_cnt >= bagel3_x+30 && h_cnt <= bagel3_x+32 && v_cnt >= bagel3_y+20 && v_cnt <= bagel3_y+24)||(h_cnt >= bagel3_x+28 && h_cnt <= bagel3_x+30 && v_cnt >= bagel3_y+22 && v_cnt <= bagel3_y+26)||(h_cnt >= bagel3_x+24 && h_cnt <= bagel3_x+28 && v_cnt >= bagel3_y+24 && v_cnt <= bagel3_y+28)||(h_cnt >= bagel3_x+14 && h_cnt <= bagel3_x+26 && v_cnt >= bagel3_y+26 && v_cnt <= bagel3_y+30)||(h_cnt >= bagel3_x+10 && h_cnt <= bagel3_x+14 && v_cnt >= bagel3_y+26 && v_cnt <= bagel3_y+28)||(h_cnt >= bagel3_x+8 && h_cnt <= bagel3_x+12 && v_cnt >= bagel3_y+24 && v_cnt <= bagel3_y+26)||(h_cnt >= bagel3_x+6 && h_cnt <= bagel3_x+12 && v_cnt >= bagel3_y+8 && v_cnt <= bagel3_y+10))
					{vgaRed, vgaGreen, vgaBlue} = 12'hf69; // light pink
				else if((h_cnt >= bagel3_x+12 && h_cnt <= bagel3_x+14 && v_cnt >= bagel3_y+2 && v_cnt <= bagel3_y+4)||(h_cnt >= bagel3_x+28 && h_cnt <= bagel3_x+30 && v_cnt >= bagel3_y+4 && v_cnt <= bagel3_y+6)||(h_cnt >= bagel3_x+30 && h_cnt <= bagel3_x+32 && v_cnt >= bagel3_y+6 && v_cnt <= bagel3_y+8)||(h_cnt >= bagel3_x+32 && h_cnt <= bagel3_x+34 && v_cnt >= bagel3_y+8 && v_cnt <= bagel3_y+10)||(h_cnt >= bagel3_x+10 && h_cnt <= bagel3_x+12 && v_cnt >= bagel3_y+20 && v_cnt <= bagel3_y+22)||(h_cnt >= bagel3_x+16 && h_cnt <= bagel3_x+18 && v_cnt >= bagel3_y+20 && v_cnt <= bagel3_y+22)||(h_cnt >= bagel3_x+22 && h_cnt <= bagel3_x+24 && v_cnt >= bagel3_y+20 && v_cnt <= bagel3_y+24)||(h_cnt >= bagel3_x+6 && h_cnt <= bagel3_x+8 && v_cnt >= bagel3_y+22 && v_cnt <= bagel3_y+24)||(h_cnt >= bagel3_x+32 && h_cnt <= bagel3_x+34 && v_cnt >= bagel3_y+24 && v_cnt <= bagel3_y+28)||(h_cnt >= bagel3_x+34 && h_cnt <= bagel3_x+36 && v_cnt >= bagel3_y+22 && v_cnt <= bagel3_y+24))
					{vgaRed, vgaGreen, vgaBlue} = 12'hf48; // dark pink
				else if((h_cnt >= bagel3_x+4 && h_cnt <= bagel3_x+6 && v_cnt >= bagel3_y+24 && v_cnt <= bagel3_y+28)||(h_cnt >= bagel3_x+6 && h_cnt <= bagel3_x+8 && v_cnt >= bagel3_y+26 && v_cnt <= bagel3_y+30)||(h_cnt >= bagel3_x+8 && h_cnt <= bagel3_x+12 && v_cnt >= bagel3_y+28 && v_cnt <= bagel3_y+32)||(h_cnt >= bagel3_x+12 && h_cnt <= bagel3_x+26 && v_cnt >= bagel3_y+30 && v_cnt <= bagel3_y+34)||(h_cnt >= bagel3_x+26 && h_cnt <= bagel3_x+30 && v_cnt >= bagel3_y+28 && v_cnt <= bagel3_y+32)||(h_cnt >= bagel3_x+30 && h_cnt <= bagel3_x+32 && v_cnt >= bagel3_y+26 && v_cnt <= bagel3_y+30)||(h_cnt >= bagel3_x+4 && h_cnt <= bagel3_x+6 && v_cnt >= bagel3_y+24 && v_cnt <= bagel3_y+28)||(h_cnt >= bagel3_x+12 && h_cnt <= bagel3_x+14 && v_cnt >= bagel3_y+22 && v_cnt <= bagel3_y+24))
					{vgaRed, vgaGreen, vgaBlue} = 12'hfd5; // yellow
				
				else if((h_cnt >= bagel4_x+12 && h_cnt <= bagel4_x+26 && v_cnt >= bagel4_y && v_cnt <= bagel4_y+2)||(h_cnt >= bagel4_x+8 && h_cnt <= bagel4_x+12 && v_cnt >= bagel4_y+2 && v_cnt <= bagel4_y+4)||(h_cnt >= bagel4_x+26 && h_cnt <= bagel4_x+30 && v_cnt >= bagel4_y+2 && v_cnt <= bagel4_y+4)||(h_cnt >= bagel4_x+6 && h_cnt <= bagel4_x+8 && v_cnt >= bagel4_y+4 && v_cnt <= bagel4_y+6)||(h_cnt >= bagel4_x+30 && h_cnt <= bagel4_x+32 && v_cnt >= bagel4_y+4 && v_cnt <= bagel4_y+6)||(h_cnt >= bagel4_x+4 && h_cnt <= bagel4_x+6 && v_cnt >= bagel4_y+6 && v_cnt <= bagel4_y+8)||(h_cnt >= bagel4_x+32 && h_cnt <= bagel4_x+34 && v_cnt >= bagel4_y+6 && v_cnt <= bagel4_y+8)||(h_cnt >= bagel4_x+2 && h_cnt <= bagel4_x+4 && v_cnt >= bagel4_y+8 && v_cnt <= bagel4_y+12)||(h_cnt >= bagel4_x+34 && h_cnt <= bagel4_x+36 && v_cnt >= bagel4_y+8 && v_cnt <= bagel4_y+12)||(h_cnt >= bagel4_x && h_cnt <= bagel4_x+2 && v_cnt >= bagel4_y+12 && v_cnt <= bagel4_y+24)||(h_cnt >= bagel4_x+36 && h_cnt <= bagel4_x+38 && v_cnt >= bagel4_y+12 && v_cnt <= bagel4_y+24)||(h_cnt >= bagel4_x+2 && h_cnt <= bagel4_x+4 && v_cnt >= bagel4_y+24 && v_cnt <= bagel4_y+28)||(h_cnt >= bagel4_x+34 && h_cnt <= bagel4_x+36 && v_cnt >= bagel4_y+24 && v_cnt <= bagel4_y+28)||(h_cnt >= bagel4_x+4 && h_cnt <= bagel4_x+6 && v_cnt >= bagel4_y+28 && v_cnt <= bagel4_y+30)||(h_cnt >= bagel4_x+32 && h_cnt <= bagel4_x+34 && v_cnt >= bagel4_y+28 && v_cnt <= bagel4_y+30)||(h_cnt >= bagel4_x+6 && h_cnt <= bagel4_x+8 && v_cnt >= bagel4_y+30 && v_cnt <= bagel4_y+32)||(h_cnt >= bagel4_x+30 && h_cnt <= bagel4_x+32 && v_cnt >= bagel4_y+30 && v_cnt <= bagel4_y+32)||(h_cnt >= bagel4_x+8 && h_cnt <= bagel4_x+12 && v_cnt >= bagel4_y+32 && v_cnt <= bagel4_y+34)||(h_cnt >= bagel4_x+26 && h_cnt <= bagel4_x+30 && v_cnt >= bagel4_y+32 && v_cnt <= bagel4_y+34)||(h_cnt >= bagel4_x+12 && h_cnt <= bagel4_x+26 && v_cnt >= bagel4_y+34 && v_cnt <= bagel4_y+36)||(h_cnt >= bagel4_x+18 && h_cnt <= bagel4_x+22 && v_cnt >= bagel4_y+14 && v_cnt <= bagel4_y+16)||(h_cnt >= bagel4_x+18 && h_cnt <= bagel4_x+22 && v_cnt >= bagel4_y+20 && v_cnt <= bagel4_y+22)||(h_cnt >= bagel4_x+16 && h_cnt <= bagel4_x+18 && v_cnt >= bagel4_y+16 && v_cnt <= bagel4_y+20)||(h_cnt >= bagel4_x+22 && h_cnt <= bagel4_x+24 && v_cnt >= bagel4_y+16 && v_cnt <= bagel4_y+20))
					{vgaRed, vgaGreen, vgaBlue} = 12'h0; // black
				else if((h_cnt >= bagel4_x+14 && h_cnt <= bagel4_x+16 && v_cnt >= bagel4_y+2 && v_cnt <= bagel4_y+4)||(h_cnt >= bagel4_x+24 && h_cnt <= bagel4_x+26 && v_cnt >= bagel4_y+2 && v_cnt <= bagel4_y+4)||(h_cnt >= bagel4_x+8 && h_cnt <= bagel4_x+10 && v_cnt >= bagel4_y+4 && v_cnt <= bagel4_y+6)||(h_cnt >= bagel4_x+26 && h_cnt <= bagel4_x+28 && v_cnt >= bagel4_y+4 && v_cnt <= bagel4_y+6)||(h_cnt >= bagel4_x+6 && h_cnt <= bagel4_x+8 && v_cnt >= bagel4_y+6 && v_cnt <= bagel4_y+8)||(h_cnt >= bagel4_x+14 && h_cnt <= bagel4_x+26 && v_cnt >= bagel4_y+6 && v_cnt <= bagel4_y+8)||(h_cnt >= bagel4_x+28 && h_cnt <= bagel4_x+30 && v_cnt >= bagel4_y+6 && v_cnt <= bagel4_y+8)||(h_cnt >= bagel4_x+4 && h_cnt <= bagel4_x+6 && v_cnt >= bagel4_y+8 && v_cnt <= bagel4_y+10)||(h_cnt >= bagel4_x+12 && h_cnt <= bagel4_x+26 && v_cnt >= bagel4_y+8 && v_cnt <= bagel4_y+10)||(h_cnt >= bagel4_x+28 && h_cnt <= bagel4_x+32 && v_cnt >= bagel4_y+8 && v_cnt <= bagel4_y+10)||(h_cnt >= bagel4_x+10 && h_cnt <= bagel4_x+14 && v_cnt >= bagel4_y+10 && v_cnt <= bagel4_y+20)||(h_cnt >= bagel4_x+24 && h_cnt <= bagel4_x+26 && v_cnt >= bagel4_y+10 && v_cnt <= bagel4_y+14)||(h_cnt >= bagel4_x+30 && h_cnt <= bagel4_x+34 && v_cnt >= bagel4_y+10 && v_cnt <= bagel4_y+18)||(h_cnt >= bagel4_x+28 && h_cnt <= bagel4_x+32 && v_cnt >= bagel4_y+18 && v_cnt <= bagel4_y+20)||(h_cnt >= bagel4_x+4 && h_cnt <= bagel4_x+6 && v_cnt >= bagel4_y+18 && v_cnt <= bagel4_y+20)||(h_cnt >= bagel4_x+6 && h_cnt <= bagel4_x+10 && v_cnt >= bagel4_y+20 && v_cnt <= bagel4_y+22)||(h_cnt >= bagel4_x+12 && h_cnt <= bagel4_x+16 && v_cnt >= bagel4_y+20 && v_cnt <= bagel4_y+22)||(h_cnt >= bagel4_x+26 && h_cnt <= bagel4_x+30 && v_cnt >= bagel4_y+20 && v_cnt <= bagel4_y+22)||(h_cnt >= bagel4_x+34 && h_cnt <= bagel4_x+36 && v_cnt >= bagel4_y+20 && v_cnt <= bagel4_y+22)||(h_cnt >= bagel4_x+4 && h_cnt <= bagel4_x+6 && v_cnt >= bagel4_y+22 && v_cnt <= bagel4_y+24)||(h_cnt >= bagel4_x+8 && h_cnt <= bagel4_x+12 && v_cnt >= bagel4_y+22 && v_cnt <= bagel4_y+24)||(h_cnt >= bagel4_x+14 && h_cnt <= bagel4_x+22 && v_cnt >= bagel4_y+22 && v_cnt <= bagel4_y+24)||(h_cnt >= bagel4_x+24 && h_cnt <= bagel4_x+28 && v_cnt >= bagel4_y+22 && v_cnt <= bagel4_y+24)||(h_cnt >= bagel4_x+32 && h_cnt <= bagel4_x+34 && v_cnt >= bagel4_y+22 && v_cnt <= bagel4_y+24)||(h_cnt >= bagel4_x+6 && h_cnt <= bagel4_x+8 && v_cnt >= bagel4_y+24 && v_cnt <= bagel4_y+26)||(h_cnt >= bagel4_x+12 && h_cnt <= bagel4_x+24 && v_cnt >= bagel4_y+24 && v_cnt <= bagel4_y+26)||(h_cnt >= bagel4_x+30 && h_cnt <= bagel4_x+32 && v_cnt >= bagel4_y+24 && v_cnt <= bagel4_y+26)||(h_cnt >= bagel4_x+8 && h_cnt <= bagel4_x+10 && v_cnt >= bagel4_y+26 && v_cnt <= bagel4_y+28)||(h_cnt >= bagel4_x+28 && h_cnt <= bagel4_x+30 && v_cnt >= bagel4_y+26 && v_cnt <= bagel4_y+28)||(h_cnt >= bagel4_x+12 && h_cnt <= bagel4_x+14 && v_cnt >= bagel4_y+28 && v_cnt <= bagel4_y+30)||(h_cnt >= bagel4_x+24 && h_cnt <= bagel4_x+26 && v_cnt >= bagel4_y+28 && v_cnt <= bagel4_y+30))
					{vgaRed, vgaGreen, vgaBlue} = 12'hf9c; // baby pink
				else if((h_cnt >= bagel4_x+16 && h_cnt <= bagel4_x+24 && v_cnt >= bagel4_y+2 && v_cnt <= bagel4_y+4)||(h_cnt >= bagel4_x+10 && h_cnt <= bagel4_x+26 && v_cnt >= bagel4_y+4 && v_cnt <= bagel4_y+6)||(h_cnt >= bagel4_x+8 && h_cnt <= bagel4_x+14 && v_cnt >= bagel4_y+6 && v_cnt <= bagel4_y+8)||(h_cnt >= bagel4_x+26 && h_cnt <= bagel4_x+28 && v_cnt >= bagel4_y+6 && v_cnt <= bagel4_y+20)||(h_cnt >= bagel4_x+28 && h_cnt <= bagel4_x+30 && v_cnt >= bagel4_y+10 && v_cnt <= bagel4_y+18)||(h_cnt >= bagel4_x+24 && h_cnt <= bagel4_x+26 && v_cnt >= bagel4_y+14 && v_cnt <= bagel4_y+22)||(h_cnt >= bagel4_x+14 && h_cnt <= bagel4_x+24 && v_cnt >= bagel4_y+10 && v_cnt <= bagel4_y+14)||(h_cnt >= bagel4_x+4 && h_cnt <= bagel4_x+10 && v_cnt >= bagel4_y+10 && v_cnt <= bagel4_y+18)||(h_cnt >= bagel4_x+2 && h_cnt <= bagel4_x+4 && v_cnt >= bagel4_y+12 && v_cnt <= bagel4_y+24)||(h_cnt >= bagel4_x+6 && h_cnt <= bagel4_x+10 && v_cnt >= bagel4_y+18 && v_cnt <= bagel4_y+20)||(h_cnt >= bagel4_x+4 && h_cnt <= bagel4_x+6 && v_cnt >= bagel4_y+20 && v_cnt <= bagel4_y+22)||(h_cnt >= bagel4_x+34 && h_cnt <= bagel4_x+36 && v_cnt >= bagel4_y+12 && v_cnt <= bagel4_y+20)||(h_cnt >= bagel4_x+22 && h_cnt <= bagel4_x+24 && v_cnt >= bagel4_y+14 && v_cnt <= bagel4_y+16)||(h_cnt >= bagel4_x+14 && h_cnt <= bagel4_x+18 && v_cnt >= bagel4_y+14 && v_cnt <= bagel4_y+16)||(h_cnt >= bagel4_x+14 && h_cnt <= bagel4_x+16 && v_cnt >= bagel4_y+16 && v_cnt <= bagel4_y+20)||(h_cnt >= bagel4_x+32 && h_cnt <= bagel4_x+34 && v_cnt >= bagel4_y+18 && v_cnt <= bagel4_y+22)||(h_cnt >= bagel4_x+30 && h_cnt <= bagel4_x+32 && v_cnt >= bagel4_y+20 && v_cnt <= bagel4_y+24)||(h_cnt >= bagel4_x+28 && h_cnt <= bagel4_x+30 && v_cnt >= bagel4_y+22 && v_cnt <= bagel4_y+26)||(h_cnt >= bagel4_x+24 && h_cnt <= bagel4_x+28 && v_cnt >= bagel4_y+24 && v_cnt <= bagel4_y+28)||(h_cnt >= bagel4_x+14 && h_cnt <= bagel4_x+26 && v_cnt >= bagel4_y+26 && v_cnt <= bagel4_y+30)||(h_cnt >= bagel4_x+10 && h_cnt <= bagel4_x+14 && v_cnt >= bagel4_y+26 && v_cnt <= bagel4_y+28)||(h_cnt >= bagel4_x+8 && h_cnt <= bagel4_x+12 && v_cnt >= bagel4_y+24 && v_cnt <= bagel4_y+26)||(h_cnt >= bagel4_x+6 && h_cnt <= bagel4_x+12 && v_cnt >= bagel4_y+8 && v_cnt <= bagel4_y+10))
					{vgaRed, vgaGreen, vgaBlue} = 12'hf69; // light pink
				else if((h_cnt >= bagel4_x+12 && h_cnt <= bagel4_x+14 && v_cnt >= bagel4_y+2 && v_cnt <= bagel4_y+4)||(h_cnt >= bagel4_x+28 && h_cnt <= bagel4_x+30 && v_cnt >= bagel4_y+4 && v_cnt <= bagel4_y+6)||(h_cnt >= bagel4_x+30 && h_cnt <= bagel4_x+32 && v_cnt >= bagel4_y+6 && v_cnt <= bagel4_y+8)||(h_cnt >= bagel4_x+32 && h_cnt <= bagel4_x+34 && v_cnt >= bagel4_y+8 && v_cnt <= bagel4_y+10)||(h_cnt >= bagel4_x+10 && h_cnt <= bagel4_x+12 && v_cnt >= bagel4_y+20 && v_cnt <= bagel4_y+22)||(h_cnt >= bagel4_x+16 && h_cnt <= bagel4_x+18 && v_cnt >= bagel4_y+20 && v_cnt <= bagel4_y+22)||(h_cnt >= bagel4_x+22 && h_cnt <= bagel4_x+24 && v_cnt >= bagel4_y+20 && v_cnt <= bagel4_y+24)||(h_cnt >= bagel4_x+6 && h_cnt <= bagel4_x+8 && v_cnt >= bagel4_y+22 && v_cnt <= bagel4_y+24)||(h_cnt >= bagel4_x+32 && h_cnt <= bagel4_x+34 && v_cnt >= bagel4_y+24 && v_cnt <= bagel4_y+28)||(h_cnt >= bagel4_x+34 && h_cnt <= bagel4_x+36 && v_cnt >= bagel4_y+22 && v_cnt <= bagel4_y+24))
					{vgaRed, vgaGreen, vgaBlue} = 12'hf48; // dark pink
				else if((h_cnt >= bagel4_x+4 && h_cnt <= bagel4_x+6 && v_cnt >= bagel4_y+24 && v_cnt <= bagel4_y+28)||(h_cnt >= bagel4_x+6 && h_cnt <= bagel4_x+8 && v_cnt >= bagel4_y+26 && v_cnt <= bagel4_y+30)||(h_cnt >= bagel4_x+8 && h_cnt <= bagel4_x+12 && v_cnt >= bagel4_y+28 && v_cnt <= bagel4_y+32)||(h_cnt >= bagel4_x+12 && h_cnt <= bagel4_x+26 && v_cnt >= bagel4_y+30 && v_cnt <= bagel4_y+34)||(h_cnt >= bagel4_x+26 && h_cnt <= bagel4_x+30 && v_cnt >= bagel4_y+28 && v_cnt <= bagel4_y+32)||(h_cnt >= bagel4_x+30 && h_cnt <= bagel4_x+32 && v_cnt >= bagel4_y+26 && v_cnt <= bagel4_y+30)||(h_cnt >= bagel4_x+4 && h_cnt <= bagel4_x+6 && v_cnt >= bagel4_y+24 && v_cnt <= bagel4_y+28)||(h_cnt >= bagel4_x+12 && h_cnt <= bagel4_x+14 && v_cnt >= bagel4_y+22 && v_cnt <= bagel4_y+24))
					{vgaRed, vgaGreen, vgaBlue} = 12'hfd5; // yellow
				
				else if((h_cnt >= bagel5_x+12 && h_cnt <= bagel5_x+26 && v_cnt >= bagel5_y && v_cnt <= bagel5_y+2)||(h_cnt >= bagel5_x+8 && h_cnt <= bagel5_x+12 && v_cnt >= bagel5_y+2 && v_cnt <= bagel5_y+4)||(h_cnt >= bagel5_x+26 && h_cnt <= bagel5_x+30 && v_cnt >= bagel5_y+2 && v_cnt <= bagel5_y+4)||(h_cnt >= bagel5_x+6 && h_cnt <= bagel5_x+8 && v_cnt >= bagel5_y+4 && v_cnt <= bagel5_y+6)||(h_cnt >= bagel5_x+30 && h_cnt <= bagel5_x+32 && v_cnt >= bagel5_y+4 && v_cnt <= bagel5_y+6)||(h_cnt >= bagel5_x+4 && h_cnt <= bagel5_x+6 && v_cnt >= bagel5_y+6 && v_cnt <= bagel5_y+8)||(h_cnt >= bagel5_x+32 && h_cnt <= bagel5_x+34 && v_cnt >= bagel5_y+6 && v_cnt <= bagel5_y+8)||(h_cnt >= bagel5_x+2 && h_cnt <= bagel5_x+4 && v_cnt >= bagel5_y+8 && v_cnt <= bagel5_y+12)||(h_cnt >= bagel5_x+34 && h_cnt <= bagel5_x+36 && v_cnt >= bagel5_y+8 && v_cnt <= bagel5_y+12)||(h_cnt >= bagel5_x && h_cnt <= bagel5_x+2 && v_cnt >= bagel5_y+12 && v_cnt <= bagel5_y+24)||(h_cnt >= bagel5_x+36 && h_cnt <= bagel5_x+38 && v_cnt >= bagel5_y+12 && v_cnt <= bagel5_y+24)||(h_cnt >= bagel5_x+2 && h_cnt <= bagel5_x+4 && v_cnt >= bagel5_y+24 && v_cnt <= bagel5_y+28)||(h_cnt >= bagel5_x+34 && h_cnt <= bagel5_x+36 && v_cnt >= bagel5_y+24 && v_cnt <= bagel5_y+28)||(h_cnt >= bagel5_x+4 && h_cnt <= bagel5_x+6 && v_cnt >= bagel5_y+28 && v_cnt <= bagel5_y+30)||(h_cnt >= bagel5_x+32 && h_cnt <= bagel5_x+34 && v_cnt >= bagel5_y+28 && v_cnt <= bagel5_y+30)||(h_cnt >= bagel5_x+6 && h_cnt <= bagel5_x+8 && v_cnt >= bagel5_y+30 && v_cnt <= bagel5_y+32)||(h_cnt >= bagel5_x+30 && h_cnt <= bagel5_x+32 && v_cnt >= bagel5_y+30 && v_cnt <= bagel5_y+32)||(h_cnt >= bagel5_x+8 && h_cnt <= bagel5_x+12 && v_cnt >= bagel5_y+32 && v_cnt <= bagel5_y+34)||(h_cnt >= bagel5_x+26 && h_cnt <= bagel5_x+30 && v_cnt >= bagel5_y+32 && v_cnt <= bagel5_y+34)||(h_cnt >= bagel5_x+12 && h_cnt <= bagel5_x+26 && v_cnt >= bagel5_y+34 && v_cnt <= bagel5_y+36)||(h_cnt >= bagel5_x+18 && h_cnt <= bagel5_x+22 && v_cnt >= bagel5_y+14 && v_cnt <= bagel5_y+16)||(h_cnt >= bagel5_x+18 && h_cnt <= bagel5_x+22 && v_cnt >= bagel5_y+20 && v_cnt <= bagel5_y+22)||(h_cnt >= bagel5_x+16 && h_cnt <= bagel5_x+18 && v_cnt >= bagel5_y+16 && v_cnt <= bagel5_y+20)||(h_cnt >= bagel5_x+22 && h_cnt <= bagel5_x+24 && v_cnt >= bagel5_y+16 && v_cnt <= bagel5_y+20))
					{vgaRed, vgaGreen, vgaBlue} = 12'h0; // black
				else if((h_cnt >= bagel5_x+14 && h_cnt <= bagel5_x+16 && v_cnt >= bagel5_y+2 && v_cnt <= bagel5_y+4)||(h_cnt >= bagel5_x+24 && h_cnt <= bagel5_x+26 && v_cnt >= bagel5_y+2 && v_cnt <= bagel5_y+4)||(h_cnt >= bagel5_x+8 && h_cnt <= bagel5_x+10 && v_cnt >= bagel5_y+4 && v_cnt <= bagel5_y+6)||(h_cnt >= bagel5_x+26 && h_cnt <= bagel5_x+28 && v_cnt >= bagel5_y+4 && v_cnt <= bagel5_y+6)||(h_cnt >= bagel5_x+6 && h_cnt <= bagel5_x+8 && v_cnt >= bagel5_y+6 && v_cnt <= bagel5_y+8)||(h_cnt >= bagel5_x+14 && h_cnt <= bagel5_x+26 && v_cnt >= bagel5_y+6 && v_cnt <= bagel5_y+8)||(h_cnt >= bagel5_x+28 && h_cnt <= bagel5_x+30 && v_cnt >= bagel5_y+6 && v_cnt <= bagel5_y+8)||(h_cnt >= bagel5_x+4 && h_cnt <= bagel5_x+6 && v_cnt >= bagel5_y+8 && v_cnt <= bagel5_y+10)||(h_cnt >= bagel5_x+12 && h_cnt <= bagel5_x+26 && v_cnt >= bagel5_y+8 && v_cnt <= bagel5_y+10)||(h_cnt >= bagel5_x+28 && h_cnt <= bagel5_x+32 && v_cnt >= bagel5_y+8 && v_cnt <= bagel5_y+10)||(h_cnt >= bagel5_x+10 && h_cnt <= bagel5_x+14 && v_cnt >= bagel5_y+10 && v_cnt <= bagel5_y+20)||(h_cnt >= bagel5_x+24 && h_cnt <= bagel5_x+26 && v_cnt >= bagel5_y+10 && v_cnt <= bagel5_y+14)||(h_cnt >= bagel5_x+30 && h_cnt <= bagel5_x+34 && v_cnt >= bagel5_y+10 && v_cnt <= bagel5_y+18)||(h_cnt >= bagel5_x+28 && h_cnt <= bagel5_x+32 && v_cnt >= bagel5_y+18 && v_cnt <= bagel5_y+20)||(h_cnt >= bagel5_x+4 && h_cnt <= bagel5_x+6 && v_cnt >= bagel5_y+18 && v_cnt <= bagel5_y+20)||(h_cnt >= bagel5_x+6 && h_cnt <= bagel5_x+10 && v_cnt >= bagel5_y+20 && v_cnt <= bagel5_y+22)||(h_cnt >= bagel5_x+12 && h_cnt <= bagel5_x+16 && v_cnt >= bagel5_y+20 && v_cnt <= bagel5_y+22)||(h_cnt >= bagel5_x+26 && h_cnt <= bagel5_x+30 && v_cnt >= bagel5_y+20 && v_cnt <= bagel5_y+22)||(h_cnt >= bagel5_x+34 && h_cnt <= bagel5_x+36 && v_cnt >= bagel5_y+20 && v_cnt <= bagel5_y+22)||(h_cnt >= bagel5_x+4 && h_cnt <= bagel5_x+6 && v_cnt >= bagel5_y+22 && v_cnt <= bagel5_y+24)||(h_cnt >= bagel5_x+8 && h_cnt <= bagel5_x+12 && v_cnt >= bagel5_y+22 && v_cnt <= bagel5_y+24)||(h_cnt >= bagel5_x+14 && h_cnt <= bagel5_x+22 && v_cnt >= bagel5_y+22 && v_cnt <= bagel5_y+24)||(h_cnt >= bagel5_x+24 && h_cnt <= bagel5_x+28 && v_cnt >= bagel5_y+22 && v_cnt <= bagel5_y+24)||(h_cnt >= bagel5_x+32 && h_cnt <= bagel5_x+34 && v_cnt >= bagel5_y+22 && v_cnt <= bagel5_y+24)||(h_cnt >= bagel5_x+6 && h_cnt <= bagel5_x+8 && v_cnt >= bagel5_y+24 && v_cnt <= bagel5_y+26)||(h_cnt >= bagel5_x+12 && h_cnt <= bagel5_x+24 && v_cnt >= bagel5_y+24 && v_cnt <= bagel5_y+26)||(h_cnt >= bagel5_x+30 && h_cnt <= bagel5_x+32 && v_cnt >= bagel5_y+24 && v_cnt <= bagel5_y+26)||(h_cnt >= bagel5_x+8 && h_cnt <= bagel5_x+10 && v_cnt >= bagel5_y+26 && v_cnt <= bagel5_y+28)||(h_cnt >= bagel5_x+28 && h_cnt <= bagel5_x+30 && v_cnt >= bagel5_y+26 && v_cnt <= bagel5_y+28)||(h_cnt >= bagel5_x+12 && h_cnt <= bagel5_x+14 && v_cnt >= bagel5_y+28 && v_cnt <= bagel5_y+30)||(h_cnt >= bagel5_x+24 && h_cnt <= bagel5_x+26 && v_cnt >= bagel5_y+28 && v_cnt <= bagel5_y+30))
					{vgaRed, vgaGreen, vgaBlue} = 12'hf9c; // baby pink
				else if((h_cnt >= bagel5_x+16 && h_cnt <= bagel5_x+24 && v_cnt >= bagel5_y+2 && v_cnt <= bagel5_y+4)||(h_cnt >= bagel5_x+10 && h_cnt <= bagel5_x+26 && v_cnt >= bagel5_y+4 && v_cnt <= bagel5_y+6)||(h_cnt >= bagel5_x+8 && h_cnt <= bagel5_x+14 && v_cnt >= bagel5_y+6 && v_cnt <= bagel5_y+8)||(h_cnt >= bagel5_x+26 && h_cnt <= bagel5_x+28 && v_cnt >= bagel5_y+6 && v_cnt <= bagel5_y+20)||(h_cnt >= bagel5_x+28 && h_cnt <= bagel5_x+30 && v_cnt >= bagel5_y+10 && v_cnt <= bagel5_y+18)||(h_cnt >= bagel5_x+24 && h_cnt <= bagel5_x+26 && v_cnt >= bagel5_y+14 && v_cnt <= bagel5_y+22)||(h_cnt >= bagel5_x+14 && h_cnt <= bagel5_x+24 && v_cnt >= bagel5_y+10 && v_cnt <= bagel5_y+14)||(h_cnt >= bagel5_x+4 && h_cnt <= bagel5_x+10 && v_cnt >= bagel5_y+10 && v_cnt <= bagel5_y+18)||(h_cnt >= bagel5_x+2 && h_cnt <= bagel5_x+4 && v_cnt >= bagel5_y+12 && v_cnt <= bagel5_y+24)||(h_cnt >= bagel5_x+6 && h_cnt <= bagel5_x+10 && v_cnt >= bagel5_y+18 && v_cnt <= bagel5_y+20)||(h_cnt >= bagel5_x+4 && h_cnt <= bagel5_x+6 && v_cnt >= bagel5_y+20 && v_cnt <= bagel5_y+22)||(h_cnt >= bagel5_x+34 && h_cnt <= bagel5_x+36 && v_cnt >= bagel5_y+12 && v_cnt <= bagel5_y+20)||(h_cnt >= bagel5_x+22 && h_cnt <= bagel5_x+24 && v_cnt >= bagel5_y+14 && v_cnt <= bagel5_y+16)||(h_cnt >= bagel5_x+14 && h_cnt <= bagel5_x+18 && v_cnt >= bagel5_y+14 && v_cnt <= bagel5_y+16)||(h_cnt >= bagel5_x+14 && h_cnt <= bagel5_x+16 && v_cnt >= bagel5_y+16 && v_cnt <= bagel5_y+20)||(h_cnt >= bagel5_x+32 && h_cnt <= bagel5_x+34 && v_cnt >= bagel5_y+18 && v_cnt <= bagel5_y+22)||(h_cnt >= bagel5_x+30 && h_cnt <= bagel5_x+32 && v_cnt >= bagel5_y+20 && v_cnt <= bagel5_y+24)||(h_cnt >= bagel5_x+28 && h_cnt <= bagel5_x+30 && v_cnt >= bagel5_y+22 && v_cnt <= bagel5_y+26)||(h_cnt >= bagel5_x+24 && h_cnt <= bagel5_x+28 && v_cnt >= bagel5_y+24 && v_cnt <= bagel5_y+28)||(h_cnt >= bagel5_x+14 && h_cnt <= bagel5_x+26 && v_cnt >= bagel5_y+26 && v_cnt <= bagel5_y+30)||(h_cnt >= bagel5_x+10 && h_cnt <= bagel5_x+14 && v_cnt >= bagel5_y+26 && v_cnt <= bagel5_y+28)||(h_cnt >= bagel5_x+8 && h_cnt <= bagel5_x+12 && v_cnt >= bagel5_y+24 && v_cnt <= bagel5_y+26)||(h_cnt >= bagel5_x+6 && h_cnt <= bagel5_x+12 && v_cnt >= bagel5_y+8 && v_cnt <= bagel5_y+10))
					{vgaRed, vgaGreen, vgaBlue} = 12'hf69; // light pink
				else if((h_cnt >= bagel5_x+12 && h_cnt <= bagel5_x+14 && v_cnt >= bagel5_y+2 && v_cnt <= bagel5_y+4)||(h_cnt >= bagel5_x+28 && h_cnt <= bagel5_x+30 && v_cnt >= bagel5_y+4 && v_cnt <= bagel5_y+6)||(h_cnt >= bagel5_x+30 && h_cnt <= bagel5_x+32 && v_cnt >= bagel5_y+6 && v_cnt <= bagel5_y+8)||(h_cnt >= bagel5_x+32 && h_cnt <= bagel5_x+34 && v_cnt >= bagel5_y+8 && v_cnt <= bagel5_y+10)||(h_cnt >= bagel5_x+10 && h_cnt <= bagel5_x+12 && v_cnt >= bagel5_y+20 && v_cnt <= bagel5_y+22)||(h_cnt >= bagel5_x+16 && h_cnt <= bagel5_x+18 && v_cnt >= bagel5_y+20 && v_cnt <= bagel5_y+22)||(h_cnt >= bagel5_x+22 && h_cnt <= bagel5_x+24 && v_cnt >= bagel5_y+20 && v_cnt <= bagel5_y+24)||(h_cnt >= bagel5_x+6 && h_cnt <= bagel5_x+8 && v_cnt >= bagel5_y+22 && v_cnt <= bagel5_y+24)||(h_cnt >= bagel5_x+32 && h_cnt <= bagel5_x+34 && v_cnt >= bagel5_y+24 && v_cnt <= bagel5_y+28)||(h_cnt >= bagel5_x+34 && h_cnt <= bagel5_x+36 && v_cnt >= bagel5_y+22 && v_cnt <= bagel5_y+24))
					{vgaRed, vgaGreen, vgaBlue} = 12'hf48; // dark pink
				else if((h_cnt >= bagel5_x+4 && h_cnt <= bagel5_x+6 && v_cnt >= bagel5_y+24 && v_cnt <= bagel5_y+28)||(h_cnt >= bagel5_x+6 && h_cnt <= bagel5_x+8 && v_cnt >= bagel5_y+26 && v_cnt <= bagel5_y+30)||(h_cnt >= bagel5_x+8 && h_cnt <= bagel5_x+12 && v_cnt >= bagel5_y+28 && v_cnt <= bagel5_y+32)||(h_cnt >= bagel5_x+12 && h_cnt <= bagel5_x+26 && v_cnt >= bagel5_y+30 && v_cnt <= bagel5_y+34)||(h_cnt >= bagel5_x+26 && h_cnt <= bagel5_x+30 && v_cnt >= bagel5_y+28 && v_cnt <= bagel5_y+32)||(h_cnt >= bagel5_x+30 && h_cnt <= bagel5_x+32 && v_cnt >= bagel5_y+26 && v_cnt <= bagel5_y+30)||(h_cnt >= bagel5_x+4 && h_cnt <= bagel5_x+6 && v_cnt >= bagel5_y+24 && v_cnt <= bagel5_y+28)||(h_cnt >= bagel5_x+12 && h_cnt <= bagel5_x+14 && v_cnt >= bagel5_y+22 && v_cnt <= bagel5_y+24))
					{vgaRed, vgaGreen, vgaBlue} = 12'hfd5; // yellowelse */
				else
					{vgaRed, vgaGreen, vgaBlue} = pixel;
			end
			3'b010:begin
				if(!valid)
					{vgaRed, vgaGreen, vgaBlue} = 12'h0;
				else if(((h_cnt>=80&&h_cnt<160)&&(v_cnt>=60&&v_cnt<80))||((h_cnt>=80&&h_cnt<100)&&(v_cnt>=80&&v_cnt<200))||((h_cnt>=120&&h_cnt<160)&&(v_cnt>=120&&v_cnt<140))||((h_cnt>=80&&h_cnt<160)&&(v_cnt>=180&&v_cnt<200))||((h_cnt>=140&&h_cnt<160)&&(v_cnt>=140&&v_cnt<180)))
					{vgaRed, vgaGreen, vgaBlue} = 12'h73a; //G
				else if(((h_cnt>=180&&h_cnt<260)&&(v_cnt>=60&&v_cnt<80))||((h_cnt>=180&&h_cnt<200)&&(v_cnt>=80&&v_cnt<200))||((h_cnt>=240&&h_cnt<260)&&(v_cnt>=80&&v_cnt<200))||((h_cnt>=200&&h_cnt<240)&&(v_cnt>=120&&v_cnt<140)))
					 {vgaRed, vgaGreen, vgaBlue} = 12'h39f;//A 
				else if(((h_cnt>=280&&h_cnt<380)&&(v_cnt>=60&&v_cnt<80))||((h_cnt>=280&&h_cnt<300)&&(v_cnt>=80&&v_cnt<200))||((h_cnt>=320&&h_cnt<340)&&(v_cnt>=80&&v_cnt<200))||((h_cnt>=360&&h_cnt<380)&&(v_cnt>=80&&v_cnt<200)))
					 {vgaRed, vgaGreen, vgaBlue} = 12'h6f6;//M
				else if(((h_cnt>=400&&h_cnt<480)&&(v_cnt>=60&&v_cnt<80))||((h_cnt>=400&&h_cnt<420)&&(v_cnt>=80&&v_cnt<200))||((h_cnt>=420&&h_cnt<480)&&(v_cnt>=120&&v_cnt<140))||((h_cnt>=420&&h_cnt<480)&&(v_cnt>=180&&v_cnt<200)))
					 {vgaRed, vgaGreen, vgaBlue} = 12'hff0;//E               
				else if(((h_cnt>=80&&h_cnt<160)&&(v_cnt>=280&&v_cnt<300))||((h_cnt>=80&&h_cnt<100)&&(v_cnt>=300&&v_cnt<420))||((h_cnt>=100&&h_cnt<160)&&(v_cnt>=400&&v_cnt<420))||((h_cnt>=140&&h_cnt<160)&&(v_cnt>=300&&v_cnt<400)))
					 {vgaRed, vgaGreen, vgaBlue} = 12'hf90;//O
				else if(((h_cnt>=180&&h_cnt<200)&&(v_cnt>=280&&v_cnt<420))||((h_cnt>=240&&h_cnt<260)&&(v_cnt>=280&&v_cnt<420))||((h_cnt>=200&&h_cnt<240)&&(v_cnt>=400&&v_cnt<420)))
					 {vgaRed, vgaGreen, vgaBlue} = 12'hf00;//V
				else if(((h_cnt>=280&&h_cnt<360)&&(v_cnt>=280&&v_cnt<300))||((h_cnt>=300&&h_cnt<360)&&(v_cnt>=340&&v_cnt<360))||((h_cnt>=300&&h_cnt<360)&&(v_cnt>=400&&v_cnt<420))||((h_cnt>=280&&h_cnt<300)&&(v_cnt>=300&&v_cnt<420)))
					 {vgaRed, vgaGreen, vgaBlue} = 12'hf9c;//E
				else if(((h_cnt>=380&&h_cnt<460)&&(v_cnt>=280&&v_cnt<300))||((h_cnt>=380&&h_cnt<400)&&(v_cnt>=300&&v_cnt<420))||((h_cnt>=440&&h_cnt<460)&&(v_cnt>=300&&v_cnt<360))||((h_cnt>=400&&h_cnt<440)&&(v_cnt>=340&&v_cnt<360))||((h_cnt>=400&&h_cnt<420)&&(v_cnt>=360&&v_cnt<380))||((h_cnt>=420&&h_cnt<440)&&(v_cnt>=380&&v_cnt<400))||((h_cnt>=440&&h_cnt<480)&&(v_cnt>=400&&v_cnt<420)))
					 {vgaRed, vgaGreen, vgaBlue} = 12'hfa2;//R
				else if(((h_cnt>=520&&h_cnt<540)&&(v_cnt>=280&&v_cnt<380))||((h_cnt>=560&&h_cnt<580)&&(v_cnt>=280&&v_cnt<380))||((h_cnt>=520&&h_cnt<540)&&(v_cnt>=400&&v_cnt<420))||((h_cnt>=560&&h_cnt<580)&&(v_cnt>=400&&v_cnt<420)))
					{vgaRed, vgaGreen, vgaBlue} = 12'hfff;//!!
				else
					 {vgaRed, vgaGreen, vgaBlue} = 12'hbde;	
			end
			
			3'b011:begin
			if(!valid)
					 {vgaRed, vgaGreen, vgaBlue} = 12'h0;
				else if(((h_cnt>=x+66&&h_cnt<x+72)&&(v_cnt>=370&&v_cnt<375))||((h_cnt>=x+54&&h_cnt<x+60)&&(v_cnt>=370&&v_cnt<380))||((h_cnt>=x+54&&h_cnt<x+78)&&(v_cnt>=390&&v_cnt<395))||((h_cnt>=x+60&&h_cnt<x+66)&&(v_cnt>=385&&v_cnt<390)))
					{vgaRed, vgaGreen, vgaBlue} = 12'h001;//BLACK
				else if(((h_cnt>=x+36&&h_cnt<x+42)&&(v_cnt>=400&&v_cnt<405))||((h_cnt>=x+60&&h_cnt<x+66)&&(v_cnt>=400&&v_cnt<405))||((h_cnt>=x+42&&h_cnt<x+48)&&(v_cnt>=405&&v_cnt<420))||((h_cnt>=x+48&&h_cnt<x+66)&&(v_cnt>=410&&v_cnt<415))||((h_cnt>=x+66&&h_cnt<x+72)&&(v_cnt>=405&&v_cnt<410))||((h_cnt>=x+72&&h_cnt<x+84)&&(v_cnt>=410&&v_cnt<425))||((h_cnt>=x+54&&h_cnt<x+72)&&(v_cnt>=415&&v_cnt<425))||((h_cnt>=x+24&&h_cnt<x+60)&&(v_cnt>=425&&v_cnt<430))||((h_cnt>=x+24&&h_cnt<x+54)&&(v_cnt>=420&&v_cnt<425))||((h_cnt>=x+24&&h_cnt<x+30)&&(v_cnt>=415&&v_cnt<420))||((h_cnt>=x+36&&h_cnt<x+42)&&(v_cnt>=415&&v_cnt<420)))
					{vgaRed, vgaGreen, vgaBlue} = 12'h00f;//BLUE
				else if(((h_cnt>=x+66&&h_cnt<x+72)&&(v_cnt>=410&&v_cnt<415))||((h_cnt>=x+48&&h_cnt<x+54)&&(v_cnt>=415&&v_cnt<420)))
					{vgaRed, vgaGreen, vgaBlue} = 12'hff0;//Y
				else if(((h_cnt>=x+90&&h_cnt<x+96)&&(v_cnt>=400&&v_cnt<425))||((h_cnt>=x+84&&h_cnt<x+90)&&(v_cnt>=405&&v_cnt<425))||((h_cnt>=x+18&&h_cnt<x+24)&&(v_cnt>=375&&v_cnt<405))||((h_cnt>=x+24&&h_cnt<x+42)&&(v_cnt>=370&&v_cnt<375))||((h_cnt>=x+30&&h_cnt<x+36)&&(v_cnt>=375&&v_cnt<390))||((h_cnt>=x+24&&h_cnt<x+30)&&(v_cnt>=390&&v_cnt<395))||((h_cnt>=x+36&&h_cnt<x+42)&&(v_cnt>=385&&v_cnt<390))||((h_cnt>=x+6&&h_cnt<x+18)&&(v_cnt>=425&&v_cnt<435))||((h_cnt>=x+12&&h_cnt<x+30)&&(v_cnt>=420&&v_cnt<425))||((h_cnt>=x+18&&h_cnt<x+24)&&(v_cnt>=425&&v_cnt<430)))
					{vgaRed, vgaGreen, vgaBlue} = 12'hfa2;              
				else if(((h_cnt>=x+72&&h_cnt<x+90)&&(v_cnt>=360&&v_cnt<365))||((h_cnt>=x+78&&h_cnt<x+90)&&(v_cnt>=365&&v_cnt<370))||((h_cnt>=x+60&&h_cnt<x+66)&&(v_cnt>=370&&v_cnt<395))||((h_cnt>=x+66&&h_cnt<x+72)&&(v_cnt>=375&&v_cnt<390))||((h_cnt>=x+72&&h_cnt<x+78)&&(v_cnt>=385&&v_cnt<390))||((h_cnt>=x+78&&h_cnt<x+84)&&(v_cnt>=385&&v_cnt<390))||((h_cnt>=x+30&&h_cnt<x+54)&&(v_cnt>=390&&v_cnt<400))||((h_cnt>=x+42&&h_cnt<x+54)&&(v_cnt>=370&&v_cnt<390))||((h_cnt>=x+24&&h_cnt<x+30)&&(v_cnt>=375&&v_cnt<390))||((h_cnt>=x+36&&h_cnt<x+42)&&(v_cnt>=375&&v_cnt<385))||((h_cnt>=x+54&&h_cnt<x+72)&&(v_cnt>=395&&v_cnt<400))||((h_cnt>=x+54&&h_cnt<x+60)&&(v_cnt>=380&&v_cnt<390))||((h_cnt>=x+0&&h_cnt<x+12)&&(v_cnt>=405&&v_cnt<415))||((h_cnt>=x+18&&h_cnt<x+24)&&(v_cnt>=410&&v_cnt<415))||((h_cnt>=x+6&&h_cnt<x+12)&&(v_cnt>=415&&v_cnt<420)))
					{vgaRed, vgaGreen, vgaBlue} = 12'hf70;
				else if(((h_cnt>=x+24&&h_cnt<x+78)&&(v_cnt>=365&&v_cnt<370))||((h_cnt>=x+30&&h_cnt<x+60)&&(v_cnt>=360&&v_cnt<365))||((h_cnt>=x+72&&h_cnt<x+90)&&(v_cnt>=370&&v_cnt<380))||((h_cnt>=x+12&&h_cnt<x+36)&&(v_cnt>=400&&v_cnt<410))||((h_cnt>=x+18&&h_cnt<x+42)&&(v_cnt>=405&&v_cnt<415))||((h_cnt>=x+42&&h_cnt<x+60)&&(v_cnt>=400&&v_cnt<405))||((h_cnt>=x+48&&h_cnt<x+66)&&(v_cnt>=405&&v_cnt<410))||((h_cnt>=x+78&&h_cnt<x+90)&&(v_cnt>=380&&v_cnt<385))||((h_cnt>=x+66&&h_cnt<x+78)&&(v_cnt>=400&&v_cnt<405))||((h_cnt>=x+72&&h_cnt<x+84)&&(v_cnt>=395&&v_cnt<400))||((h_cnt>=x+78&&h_cnt<x+84)&&(v_cnt>=390&&v_cnt<395))||((h_cnt>=x+30&&h_cnt<x+36)&&(v_cnt>=415&&v_cnt<420))||((h_cnt>=x+84&&h_cnt<x+90)&&(v_cnt>=385&&v_cnt<390)))
					{vgaRed, vgaGreen, vgaBlue} = 12'hf00;//red

				else if((h_cnt>=branch1_x+10 && h_cnt<branch1_x+12)&&(v_cnt>=branch1_y+8 && v_cnt<branch1_y+39) || (h_cnt>=branch1_x+7 && h_cnt<branch1_x+10 && v_cnt==branch1_y+10) || (h_cnt==branch1_x+6 && v_cnt>=branch1_y+8 && v_cnt<branch1_y+10) || (h_cnt==branch1_x+5 && v_cnt==branch1_y+8) || (h_cnt>=branch1_x+3 && h_cnt<branch1_x+5 && v_cnt==branch1_y+7) || (h_cnt==branch1_x+6 && v_cnt>=branch1_y+8 && v_cnt<branch1_y+10) || (h_cnt==branch1_x+2 && v_cnt>=branch1_y+5 && v_cnt<branch1_y+7) || (h_cnt==branch1_x+1 && v_cnt==branch1_y+5) || (h_cnt==branch1_x && v_cnt==branch1_y+4) || (h_cnt>=branch1_x+11 && h_cnt<branch1_x+14 && v_cnt==branch1_y+7) || (h_cnt>=branch1_x+14 && h_cnt<branch1_x+16 && v_cnt==branch1_y+5) || (h_cnt==branch1_x+14 && v_cnt==branch1_y+6) || (h_cnt>=branch1_x+16 && h_cnt<branch1_x+17 && v_cnt==branch1_y+4) || (h_cnt>=branch1_x+18 && h_cnt<branch1_x+19 && v_cnt==branch1_y+1) || (h_cnt==branch1_x+17 && v_cnt==branch1_y+3) || (h_cnt==branch1_x+18 && v_cnt==branch1_y+2))
					{vgaRed, vgaGreen, vgaBlue} = 12'h644; // brown
				else if((h_cnt>=branch1_x+5 && h_cnt<branch1_x+6 && v_cnt==branch1_y+10) || (h_cnt>=branch1_x+2 && h_cnt<branch1_x+4 && v_cnt==branch1_y+8) || (h_cnt>=branch1_x && h_cnt<branch1_x+1 && v_cnt==branch1_y+6) || (h_cnt>=branch1_x+3 && h_cnt<branch1_x+5 && v_cnt==branch1_y+6) || (h_cnt>=branch1_x+1 && h_cnt<branch1_x+2 && v_cnt==branch1_y+4) || (h_cnt>=branch1_x+13 && h_cnt<branch1_x+14 && v_cnt==branch1_y+4) || (h_cnt>=branch1_x+15 && h_cnt<branch1_x+16 && v_cnt==branch1_y+3) || (h_cnt>=branch1_x+16 && h_cnt<branch1_x+17 && v_cnt==branch1_y+5) || (h_cnt>=branch1_x+19 && h_cnt<branch1_x+20 && v_cnt==branch1_y) || (h_cnt==branch1_x+7 && v_cnt>=branch1_y+7 && v_cnt<branch1_y+8) || (h_cnt==branch1_x+17 && v_cnt>=branch1_y+1 && v_cnt<branch1_y+2) || (h_cnt==branch1_x+18 && v_cnt>=branch1_y+3 && v_cnt<branch1_y+4) || (h_cnt==branch1_x+2 && v_cnt==branch1_y+3) || (h_cnt==branch1_x+2 && v_cnt==branch1_y+7) || (h_cnt==branch1_x+4 && v_cnt==branch1_y+9) || (h_cnt==branch1_x+6 && v_cnt==branch1_y+11) || (h_cnt==branch1_x+12 && v_cnt==branch1_y+6) || (h_cnt==branch1_x+14 && v_cnt==branch1_y+8) || (h_cnt==branch1_x+19 && v_cnt==branch1_y+2) || (h_cnt==branch1_x+20 && v_cnt==branch1_y+1))
					{vgaRed, vgaGreen, vgaBlue} = 12'h9b2; // green

				else if((h_cnt>=branch2_x+10 && h_cnt<branch2_x+12)&&(v_cnt>=branch2_y+8 && v_cnt<branch2_y+39) || (h_cnt>=branch2_x+7 && h_cnt<branch2_x+10 && v_cnt==branch2_y+10) || (h_cnt==branch2_x+6 && v_cnt>=branch2_y+8 && v_cnt<branch2_y+10) || (h_cnt==branch2_x+5 && v_cnt==branch2_y+8) || (h_cnt>=branch2_x+3 && h_cnt<branch2_x+5 && v_cnt==branch2_y+7) || (h_cnt==branch2_x+6 && v_cnt>=branch2_y+8 && v_cnt<branch2_y+10) || (h_cnt==branch2_x+2 && v_cnt>=branch2_y+5 && v_cnt<branch2_y+7) || (h_cnt==branch2_x+1 && v_cnt==branch2_y+5) || (h_cnt==branch2_x && v_cnt==branch2_y+4) || (h_cnt>=branch2_x+11 && h_cnt<branch2_x+14 && v_cnt==branch2_y+7) || (h_cnt>=branch2_x+14 && h_cnt<branch2_x+16 && v_cnt==branch2_y+5) || (h_cnt==branch2_x+14 && v_cnt==branch2_y+6) || (h_cnt>=branch2_x+16 && h_cnt<branch2_x+17 && v_cnt==branch2_y+4) || (h_cnt>=branch2_x+18 && h_cnt<branch2_x+19 && v_cnt==branch2_y+1) || (h_cnt==branch2_x+17 && v_cnt==branch2_y+3) || (h_cnt==branch2_x+18 && v_cnt==branch2_y+2))
					{vgaRed, vgaGreen, vgaBlue} = 12'h644; // brown
				else if((h_cnt>=branch2_x+5 && h_cnt<branch2_x+6 && v_cnt==branch2_y+10) || (h_cnt>=branch2_x+2 && h_cnt<branch2_x+4 && v_cnt==branch2_y+8) || (h_cnt>=branch2_x && h_cnt<branch2_x+1 && v_cnt==branch2_y+6) || (h_cnt>=branch2_x+3 && h_cnt<branch2_x+5 && v_cnt==branch2_y+6) || (h_cnt>=branch2_x+1 && h_cnt<branch2_x+2 && v_cnt==branch2_y+4) || (h_cnt>=branch2_x+13 && h_cnt<branch2_x+14 && v_cnt==branch2_y+4) || (h_cnt>=branch2_x+15 && h_cnt<branch2_x+16 && v_cnt==branch2_y+3) || (h_cnt>=branch2_x+16 && h_cnt<branch2_x+17 && v_cnt==branch2_y+5) || (h_cnt>=branch2_x+19 && h_cnt<branch2_x+20 && v_cnt==branch2_y) || (h_cnt==branch2_x+7 && v_cnt>=branch2_y+7 && v_cnt<branch2_y+8) || (h_cnt==branch2_x+17 && v_cnt>=branch2_y+1 && v_cnt<branch2_y+2) || (h_cnt==branch2_x+18 && v_cnt>=branch2_y+3 && v_cnt<branch2_y+4) || (h_cnt==branch2_x+2 && v_cnt==branch2_y+3) || (h_cnt==branch2_x+2 && v_cnt==branch2_y+7) || (h_cnt==branch2_x+4 && v_cnt==branch2_y+9) || (h_cnt==branch2_x+6 && v_cnt==branch2_y+11) || (h_cnt==branch2_x+12 && v_cnt==branch2_y+6) || (h_cnt==branch2_x+14 && v_cnt==branch2_y+8) || (h_cnt==branch2_x+19 && v_cnt==branch2_y+2) || (h_cnt==branch2_x+20 && v_cnt==branch2_y+1))
					{vgaRed, vgaGreen, vgaBlue} = 12'h9b2; // green

				else if((h_cnt>=branch3_x+10 && h_cnt<branch3_x+12)&&(v_cnt>=branch3_y+8 && v_cnt<branch3_y+39) || (h_cnt>=branch3_x+7 && h_cnt<branch3_x+10 && v_cnt==branch3_y+10) || (h_cnt==branch3_x+6 && v_cnt>=branch3_y+8 && v_cnt<branch3_y+10) || (h_cnt==branch3_x+5 && v_cnt==branch3_y+8) || (h_cnt>=branch3_x+3 && h_cnt<branch3_x+5 && v_cnt==branch3_y+7) || (h_cnt==branch3_x+6 && v_cnt>=branch3_y+8 && v_cnt<branch3_y+10) || (h_cnt==branch3_x+2 && v_cnt>=branch3_y+5 && v_cnt<branch3_y+7) || (h_cnt==branch3_x+1 && v_cnt==branch3_y+5) || (h_cnt==branch3_x && v_cnt==branch3_y+4) || (h_cnt>=branch3_x+11 && h_cnt<branch3_x+14 && v_cnt==branch3_y+7) || (h_cnt>=branch3_x+14 && h_cnt<branch3_x+16 && v_cnt==branch3_y+5) || (h_cnt==branch3_x+14 && v_cnt==branch3_y+6) || (h_cnt>=branch3_x+16 && h_cnt<branch3_x+17 && v_cnt==branch3_y+4) || (h_cnt>=branch3_x+18 && h_cnt<branch3_x+19 && v_cnt==branch3_y+1) || (h_cnt==branch3_x+17 && v_cnt==branch3_y+3) || (h_cnt==branch3_x+18 && v_cnt==branch3_y+2))
					{vgaRed, vgaGreen, vgaBlue} = 12'h644; // brown
				else if((h_cnt>=branch3_x+5 && h_cnt<branch3_x+6 && v_cnt==branch3_y+10) || (h_cnt>=branch3_x+2 && h_cnt<branch3_x+4 && v_cnt==branch3_y+8) || (h_cnt>=branch3_x && h_cnt<branch3_x+1 && v_cnt==branch3_y+6) || (h_cnt>=branch3_x+3 && h_cnt<branch3_x+5 && v_cnt==branch3_y+6) || (h_cnt>=branch3_x+1 && h_cnt<branch3_x+2 && v_cnt==branch3_y+4) || (h_cnt>=branch3_x+13 && h_cnt<branch3_x+14 && v_cnt==branch3_y+4) || (h_cnt>=branch3_x+15 && h_cnt<branch3_x+16 && v_cnt==branch3_y+3) || (h_cnt>=branch3_x+16 && h_cnt<branch3_x+17 && v_cnt==branch3_y+5) || (h_cnt>=branch3_x+19 && h_cnt<branch3_x+20 && v_cnt==branch3_y) || (h_cnt==branch3_x+7 && v_cnt>=branch3_y+7 && v_cnt<branch3_y+8) || (h_cnt==branch3_x+17 && v_cnt>=branch3_y+1 && v_cnt<branch3_y+2) || (h_cnt==branch3_x+18 && v_cnt>=branch3_y+3 && v_cnt<branch3_y+4) || (h_cnt==branch3_x+2 && v_cnt==branch3_y+3) || (h_cnt==branch3_x+2 && v_cnt==branch3_y+7) || (h_cnt==branch3_x+4 && v_cnt==branch3_y+9) || (h_cnt==branch3_x+6 && v_cnt==branch3_y+11) || (h_cnt==branch3_x+12 && v_cnt==branch3_y+6) || (h_cnt==branch3_x+14 && v_cnt==branch3_y+8) || (h_cnt==branch3_x+19 && v_cnt==branch3_y+2) || (h_cnt==branch3_x+20 && v_cnt==branch3_y+1))
					{vgaRed, vgaGreen, vgaBlue} = 12'h9b2; // green

				else if((h_cnt>=branch4_x+10 && h_cnt<branch4_x+12)&&(v_cnt>=branch4_y+8 && v_cnt<branch4_y+39) || (h_cnt>=branch4_x+7 && h_cnt<branch4_x+10 && v_cnt==branch4_y+10) || (h_cnt==branch4_x+6 && v_cnt>=branch4_y+8 && v_cnt<branch4_y+10) || (h_cnt==branch4_x+5 && v_cnt==branch4_y+8) || (h_cnt>=branch4_x+3 && h_cnt<branch4_x+5 && v_cnt==branch4_y+7) || (h_cnt==branch4_x+6 && v_cnt>=branch4_y+8 && v_cnt<branch4_y+10) || (h_cnt==branch4_x+2 && v_cnt>=branch4_y+5 && v_cnt<branch4_y+7) || (h_cnt==branch4_x+1 && v_cnt==branch4_y+5) || (h_cnt==branch4_x && v_cnt==branch4_y+4) || (h_cnt>=branch4_x+11 && h_cnt<branch4_x+14 && v_cnt==branch4_y+7) || (h_cnt>=branch4_x+14 && h_cnt<branch4_x+16 && v_cnt==branch4_y+5) || (h_cnt==branch4_x+14 && v_cnt==branch4_y+6) || (h_cnt>=branch4_x+16 && h_cnt<branch4_x+17 && v_cnt==branch4_y+4) || (h_cnt>=branch4_x+18 && h_cnt<branch4_x+19 && v_cnt==branch4_y+1) || (h_cnt==branch4_x+17 && v_cnt==branch4_y+3) || (h_cnt==branch4_x+18 && v_cnt==branch4_y+2))
					{vgaRed, vgaGreen, vgaBlue} = 12'h644; // brown
				else if((h_cnt>=branch4_x+5 && h_cnt<branch4_x+6 && v_cnt==branch4_y+10) || (h_cnt>=branch4_x+2 && h_cnt<branch4_x+4 && v_cnt==branch4_y+8) || (h_cnt>=branch4_x && h_cnt<branch4_x+1 && v_cnt==branch4_y+6) || (h_cnt>=branch4_x+3 && h_cnt<branch4_x+5 && v_cnt==branch4_y+6) || (h_cnt>=branch4_x+1 && h_cnt<branch4_x+2 && v_cnt==branch4_y+4) || (h_cnt>=branch4_x+13 && h_cnt<branch4_x+14 && v_cnt==branch4_y+4) || (h_cnt>=branch4_x+15 && h_cnt<branch4_x+16 && v_cnt==branch4_y+3) || (h_cnt>=branch4_x+16 && h_cnt<branch4_x+17 && v_cnt==branch4_y+5) || (h_cnt>=branch4_x+19 && h_cnt<branch4_x+20 && v_cnt==branch4_y) || (h_cnt==branch4_x+7 && v_cnt>=branch4_y+7 && v_cnt<branch4_y+8) || (h_cnt==branch4_x+17 && v_cnt>=branch4_y+1 && v_cnt<branch4_y+2) || (h_cnt==branch4_x+18 && v_cnt>=branch4_y+3 && v_cnt<branch4_y+4) || (h_cnt==branch4_x+2 && v_cnt==branch4_y+3) || (h_cnt==branch4_x+2 && v_cnt==branch4_y+7) || (h_cnt==branch4_x+4 && v_cnt==branch4_y+9) || (h_cnt==branch4_x+6 && v_cnt==branch4_y+11) || (h_cnt==branch4_x+12 && v_cnt==branch4_y+6) || (h_cnt==branch4_x+14 && v_cnt==branch4_y+8) || (h_cnt==branch4_x+19 && v_cnt==branch4_y+2) || (h_cnt==branch4_x+20 && v_cnt==branch4_y+1))
					{vgaRed, vgaGreen, vgaBlue} = 12'h9b2; // green
					
				else if((h_cnt>=branch5_x+10 && h_cnt<branch5_x+12)&&(v_cnt>=branch5_y+8 && v_cnt<branch5_y+39) || (h_cnt>=branch5_x+7 && h_cnt<branch5_x+10 && v_cnt==branch5_y+10) || (h_cnt==branch5_x+6 && v_cnt>=branch5_y+8 && v_cnt<branch5_y+10) || (h_cnt==branch5_x+5 && v_cnt==branch5_y+8) || (h_cnt>=branch5_x+3 && h_cnt<branch5_x+5 && v_cnt==branch5_y+7) || (h_cnt==branch5_x+6 && v_cnt>=branch5_y+8 && v_cnt<branch5_y+10) || (h_cnt==branch5_x+2 && v_cnt>=branch5_y+5 && v_cnt<branch5_y+7) || (h_cnt==branch5_x+1 && v_cnt==branch5_y+5) || (h_cnt==branch5_x && v_cnt==branch5_y+4) || (h_cnt>=branch5_x+11 && h_cnt<branch5_x+14 && v_cnt==branch5_y+7) || (h_cnt>=branch5_x+14 && h_cnt<branch5_x+16 && v_cnt==branch5_y+5) || (h_cnt==branch5_x+14 && v_cnt==branch5_y+6) || (h_cnt>=branch5_x+16 && h_cnt<branch5_x+17 && v_cnt==branch5_y+4) || (h_cnt>=branch5_x+18 && h_cnt<branch5_x+19 && v_cnt==branch5_y+1) || (h_cnt==branch5_x+17 && v_cnt==branch5_y+3) || (h_cnt==branch5_x+18 && v_cnt==branch5_y+2))
					{vgaRed, vgaGreen, vgaBlue} = 12'h644; // brown
				else if((h_cnt>=branch5_x+5 && h_cnt<branch5_x+6 && v_cnt==branch5_y+10) || (h_cnt>=branch5_x+2 && h_cnt<branch5_x+4 && v_cnt==branch5_y+8) || (h_cnt>=branch5_x && h_cnt<branch5_x+1 && v_cnt==branch5_y+6) || (h_cnt>=branch5_x+3 && h_cnt<branch5_x+5 && v_cnt==branch5_y+6) || (h_cnt>=branch5_x+1 && h_cnt<branch5_x+2 && v_cnt==branch5_y+4) || (h_cnt>=branch5_x+13 && h_cnt<branch5_x+14 && v_cnt==branch5_y+4) || (h_cnt>=branch5_x+15 && h_cnt<branch5_x+16 && v_cnt==branch5_y+3) || (h_cnt>=branch5_x+16 && h_cnt<branch5_x+17 && v_cnt==branch5_y+5) || (h_cnt>=branch5_x+19 && h_cnt<branch5_x+20 && v_cnt==branch5_y) || (h_cnt==branch5_x+7 && v_cnt>=branch5_y+7 && v_cnt<branch5_y+8) || (h_cnt==branch5_x+17 && v_cnt>=branch5_y+1 && v_cnt<branch5_y+2) || (h_cnt==branch5_x+18 && v_cnt>=branch5_y+3 && v_cnt<branch5_y+4) || (h_cnt==branch5_x+2 && v_cnt==branch5_y+3) || (h_cnt==branch5_x+2 && v_cnt==branch5_y+7) || (h_cnt==branch5_x+4 && v_cnt==branch5_y+9) || (h_cnt==branch5_x+6 && v_cnt==branch5_y+11) || (h_cnt==branch5_x+12 && v_cnt==branch5_y+6) || (h_cnt==branch5_x+14 && v_cnt==branch5_y+8) || (h_cnt==branch5_x+19 && v_cnt==branch5_y+2) || (h_cnt==branch5_x+20 && v_cnt==branch5_y+1))
					{vgaRed, vgaGreen, vgaBlue} = 12'h9b2; // green
		
				else if((h_cnt >= bagel1_x+12 && h_cnt <= bagel1_x+26 && v_cnt >= bagel1_y && v_cnt <= bagel1_y+2)||(h_cnt >= bagel1_x+8 && h_cnt <= bagel1_x+12 && v_cnt >= bagel1_y+2 && v_cnt <= bagel1_y+4)||(h_cnt >= bagel1_x+26 && h_cnt <= bagel1_x+30 && v_cnt >= bagel1_y+2 && v_cnt <= bagel1_y+4)||(h_cnt >= bagel1_x+6 && h_cnt <= bagel1_x+8 && v_cnt >= bagel1_y+4 && v_cnt <= bagel1_y+6)||(h_cnt >= bagel1_x+30 && h_cnt <= bagel1_x+32 && v_cnt >= bagel1_y+4 && v_cnt <= bagel1_y+6)||(h_cnt >= bagel1_x+4 && h_cnt <= bagel1_x+6 && v_cnt >= bagel1_y+6 && v_cnt <= bagel1_y+8)||(h_cnt >= bagel1_x+32 && h_cnt <= bagel1_x+34 && v_cnt >= bagel1_y+6 && v_cnt <= bagel1_y+8)||(h_cnt >= bagel1_x+2 && h_cnt <= bagel1_x+4 && v_cnt >= bagel1_y+8 && v_cnt <= bagel1_y+12)||(h_cnt >= bagel1_x+34 && h_cnt <= bagel1_x+36 && v_cnt >= bagel1_y+8 && v_cnt <= bagel1_y+12)||(h_cnt >= bagel1_x && h_cnt <= bagel1_x+2 && v_cnt >= bagel1_y+12 && v_cnt <= bagel1_y+24)||(h_cnt >= bagel1_x+36 && h_cnt <= bagel1_x+38 && v_cnt >= bagel1_y+12 && v_cnt <= bagel1_y+24)||(h_cnt >= bagel1_x+2 && h_cnt <= bagel1_x+4 && v_cnt >= bagel1_y+24 && v_cnt <= bagel1_y+28)||(h_cnt >= bagel1_x+34 && h_cnt <= bagel1_x+36 && v_cnt >= bagel1_y+24 && v_cnt <= bagel1_y+28)||(h_cnt >= bagel1_x+4 && h_cnt <= bagel1_x+6 && v_cnt >= bagel1_y+28 && v_cnt <= bagel1_y+30)||(h_cnt >= bagel1_x+32 && h_cnt <= bagel1_x+34 && v_cnt >= bagel1_y+28 && v_cnt <= bagel1_y+30)||(h_cnt >= bagel1_x+6 && h_cnt <= bagel1_x+8 && v_cnt >= bagel1_y+30 && v_cnt <= bagel1_y+32)||(h_cnt >= bagel1_x+30 && h_cnt <= bagel1_x+32 && v_cnt >= bagel1_y+30 && v_cnt <= bagel1_y+32)||(h_cnt >= bagel1_x+8 && h_cnt <= bagel1_x+12 && v_cnt >= bagel1_y+32 && v_cnt <= bagel1_y+34)||(h_cnt >= bagel1_x+26 && h_cnt <= bagel1_x+30 && v_cnt >= bagel1_y+32 && v_cnt <= bagel1_y+34)||(h_cnt >= bagel1_x+12 && h_cnt <= bagel1_x+26 && v_cnt >= bagel1_y+34 && v_cnt <= bagel1_y+36)||(h_cnt >= bagel1_x+18 && h_cnt <= bagel1_x+22 && v_cnt >= bagel1_y+14 && v_cnt <= bagel1_y+16)||(h_cnt >= bagel1_x+18 && h_cnt <= bagel1_x+22 && v_cnt >= bagel1_y+20 && v_cnt <= bagel1_y+22)||(h_cnt >= bagel1_x+16 && h_cnt <= bagel1_x+18 && v_cnt >= bagel1_y+16 && v_cnt <= bagel1_y+20)||(h_cnt >= bagel1_x+22 && h_cnt <= bagel1_x+24 && v_cnt >= bagel1_y+16 && v_cnt <= bagel1_y+20))
					{vgaRed, vgaGreen, vgaBlue} = 12'h0; // black
				else if((h_cnt >= bagel1_x+14 && h_cnt <= bagel1_x+16 && v_cnt >= bagel1_y+2 && v_cnt <= bagel1_y+4)||(h_cnt >= bagel1_x+24 && h_cnt <= bagel1_x+26 && v_cnt >= bagel1_y+2 && v_cnt <= bagel1_y+4)||(h_cnt >= bagel1_x+8 && h_cnt <= bagel1_x+10 && v_cnt >= bagel1_y+4 && v_cnt <= bagel1_y+6)||(h_cnt >= bagel1_x+26 && h_cnt <= bagel1_x+28 && v_cnt >= bagel1_y+4 && v_cnt <= bagel1_y+6)||(h_cnt >= bagel1_x+6 && h_cnt <= bagel1_x+8 && v_cnt >= bagel1_y+6 && v_cnt <= bagel1_y+8)||(h_cnt >= bagel1_x+14 && h_cnt <= bagel1_x+26 && v_cnt >= bagel1_y+6 && v_cnt <= bagel1_y+8)||(h_cnt >= bagel1_x+28 && h_cnt <= bagel1_x+30 && v_cnt >= bagel1_y+6 && v_cnt <= bagel1_y+8)||(h_cnt >= bagel1_x+4 && h_cnt <= bagel1_x+6 && v_cnt >= bagel1_y+8 && v_cnt <= bagel1_y+10)||(h_cnt >= bagel1_x+12 && h_cnt <= bagel1_x+26 && v_cnt >= bagel1_y+8 && v_cnt <= bagel1_y+10)||(h_cnt >= bagel1_x+28 && h_cnt <= bagel1_x+32 && v_cnt >= bagel1_y+8 && v_cnt <= bagel1_y+10)||(h_cnt >= bagel1_x+10 && h_cnt <= bagel1_x+14 && v_cnt >= bagel1_y+10 && v_cnt <= bagel1_y+20)||(h_cnt >= bagel1_x+24 && h_cnt <= bagel1_x+26 && v_cnt >= bagel1_y+10 && v_cnt <= bagel1_y+14)||(h_cnt >= bagel1_x+30 && h_cnt <= bagel1_x+34 && v_cnt >= bagel1_y+10 && v_cnt <= bagel1_y+18)||(h_cnt >= bagel1_x+28 && h_cnt <= bagel1_x+32 && v_cnt >= bagel1_y+18 && v_cnt <= bagel1_y+20)||(h_cnt >= bagel1_x+4 && h_cnt <= bagel1_x+6 && v_cnt >= bagel1_y+18 && v_cnt <= bagel1_y+20)||(h_cnt >= bagel1_x+6 && h_cnt <= bagel1_x+10 && v_cnt >= bagel1_y+20 && v_cnt <= bagel1_y+22)||(h_cnt >= bagel1_x+12 && h_cnt <= bagel1_x+16 && v_cnt >= bagel1_y+20 && v_cnt <= bagel1_y+22)||(h_cnt >= bagel1_x+26 && h_cnt <= bagel1_x+30 && v_cnt >= bagel1_y+20 && v_cnt <= bagel1_y+22)||(h_cnt >= bagel1_x+34 && h_cnt <= bagel1_x+36 && v_cnt >= bagel1_y+20 && v_cnt <= bagel1_y+22)||(h_cnt >= bagel1_x+4 && h_cnt <= bagel1_x+6 && v_cnt >= bagel1_y+22 && v_cnt <= bagel1_y+24)||(h_cnt >= bagel1_x+8 && h_cnt <= bagel1_x+12 && v_cnt >= bagel1_y+22 && v_cnt <= bagel1_y+24)||(h_cnt >= bagel1_x+14 && h_cnt <= bagel1_x+22 && v_cnt >= bagel1_y+22 && v_cnt <= bagel1_y+24)||(h_cnt >= bagel1_x+24 && h_cnt <= bagel1_x+28 && v_cnt >= bagel1_y+22 && v_cnt <= bagel1_y+24)||(h_cnt >= bagel1_x+32 && h_cnt <= bagel1_x+34 && v_cnt >= bagel1_y+22 && v_cnt <= bagel1_y+24)||(h_cnt >= bagel1_x+6 && h_cnt <= bagel1_x+8 && v_cnt >= bagel1_y+24 && v_cnt <= bagel1_y+26)||(h_cnt >= bagel1_x+12 && h_cnt <= bagel1_x+24 && v_cnt >= bagel1_y+24 && v_cnt <= bagel1_y+26)||(h_cnt >= bagel1_x+30 && h_cnt <= bagel1_x+32 && v_cnt >= bagel1_y+24 && v_cnt <= bagel1_y+26)||(h_cnt >= bagel1_x+8 && h_cnt <= bagel1_x+10 && v_cnt >= bagel1_y+26 && v_cnt <= bagel1_y+28)||(h_cnt >= bagel1_x+28 && h_cnt <= bagel1_x+30 && v_cnt >= bagel1_y+26 && v_cnt <= bagel1_y+28)||(h_cnt >= bagel1_x+12 && h_cnt <= bagel1_x+14 && v_cnt >= bagel1_y+28 && v_cnt <= bagel1_y+30)||(h_cnt >= bagel1_x+24 && h_cnt <= bagel1_x+26 && v_cnt >= bagel1_y+28 && v_cnt <= bagel1_y+30))
					{vgaRed, vgaGreen, vgaBlue} = 12'hf9c; // baby pink
				else if((h_cnt >= bagel1_x+16 && h_cnt <= bagel1_x+24 && v_cnt >= bagel1_y+2 && v_cnt <= bagel1_y+4)||(h_cnt >= bagel1_x+10 && h_cnt <= bagel1_x+26 && v_cnt >= bagel1_y+4 && v_cnt <= bagel1_y+6)||(h_cnt >= bagel1_x+8 && h_cnt <= bagel1_x+14 && v_cnt >= bagel1_y+6 && v_cnt <= bagel1_y+8)||(h_cnt >= bagel1_x+26 && h_cnt <= bagel1_x+28 && v_cnt >= bagel1_y+6 && v_cnt <= bagel1_y+20)||(h_cnt >= bagel1_x+28 && h_cnt <= bagel1_x+30 && v_cnt >= bagel1_y+10 && v_cnt <= bagel1_y+18)||(h_cnt >= bagel1_x+24 && h_cnt <= bagel1_x+26 && v_cnt >= bagel1_y+14 && v_cnt <= bagel1_y+22)||(h_cnt >= bagel1_x+14 && h_cnt <= bagel1_x+24 && v_cnt >= bagel1_y+10 && v_cnt <= bagel1_y+14)||(h_cnt >= bagel1_x+4 && h_cnt <= bagel1_x+10 && v_cnt >= bagel1_y+10 && v_cnt <= bagel1_y+18)||(h_cnt >= bagel1_x+2 && h_cnt <= bagel1_x+4 && v_cnt >= bagel1_y+12 && v_cnt <= bagel1_y+24)||(h_cnt >= bagel1_x+6 && h_cnt <= bagel1_x+10 && v_cnt >= bagel1_y+18 && v_cnt <= bagel1_y+20)||(h_cnt >= bagel1_x+4 && h_cnt <= bagel1_x+6 && v_cnt >= bagel1_y+20 && v_cnt <= bagel1_y+22)||(h_cnt >= bagel1_x+34 && h_cnt <= bagel1_x+36 && v_cnt >= bagel1_y+12 && v_cnt <= bagel1_y+20)||(h_cnt >= bagel1_x+22 && h_cnt <= bagel1_x+24 && v_cnt >= bagel1_y+14 && v_cnt <= bagel1_y+16)||(h_cnt >= bagel1_x+14 && h_cnt <= bagel1_x+18 && v_cnt >= bagel1_y+14 && v_cnt <= bagel1_y+16)||(h_cnt >= bagel1_x+14 && h_cnt <= bagel1_x+16 && v_cnt >= bagel1_y+16 && v_cnt <= bagel1_y+20)||(h_cnt >= bagel1_x+32 && h_cnt <= bagel1_x+34 && v_cnt >= bagel1_y+18 && v_cnt <= bagel1_y+22)||(h_cnt >= bagel1_x+30 && h_cnt <= bagel1_x+32 && v_cnt >= bagel1_y+20 && v_cnt <= bagel1_y+24)||(h_cnt >= bagel1_x+28 && h_cnt <= bagel1_x+30 && v_cnt >= bagel1_y+22 && v_cnt <= bagel1_y+26)||(h_cnt >= bagel1_x+24 && h_cnt <= bagel1_x+28 && v_cnt >= bagel1_y+24 && v_cnt <= bagel1_y+28)||(h_cnt >= bagel1_x+14 && h_cnt <= bagel1_x+26 && v_cnt >= bagel1_y+26 && v_cnt <= bagel1_y+30)||(h_cnt >= bagel1_x+10 && h_cnt <= bagel1_x+14 && v_cnt >= bagel1_y+26 && v_cnt <= bagel1_y+28)||(h_cnt >= bagel1_x+8 && h_cnt <= bagel1_x+12 && v_cnt >= bagel1_y+24 && v_cnt <= bagel1_y+26)||(h_cnt >= bagel1_x+6 && h_cnt <= bagel1_x+12 && v_cnt >= bagel1_y+8 && v_cnt <= bagel1_y+10))
					{vgaRed, vgaGreen, vgaBlue} = 12'hf69; // light pink
				else if((h_cnt >= bagel1_x+12 && h_cnt <= bagel1_x+14 && v_cnt >= bagel1_y+2 && v_cnt <= bagel1_y+4)||(h_cnt >= bagel1_x+28 && h_cnt <= bagel1_x+30 && v_cnt >= bagel1_y+4 && v_cnt <= bagel1_y+6)||(h_cnt >= bagel1_x+30 && h_cnt <= bagel1_x+32 && v_cnt >= bagel1_y+6 && v_cnt <= bagel1_y+8)||(h_cnt >= bagel1_x+32 && h_cnt <= bagel1_x+34 && v_cnt >= bagel1_y+8 && v_cnt <= bagel1_y+10)||(h_cnt >= bagel1_x+10 && h_cnt <= bagel1_x+12 && v_cnt >= bagel1_y+20 && v_cnt <= bagel1_y+22)||(h_cnt >= bagel1_x+16 && h_cnt <= bagel1_x+18 && v_cnt >= bagel1_y+20 && v_cnt <= bagel1_y+22)||(h_cnt >= bagel1_x+22 && h_cnt <= bagel1_x+24 && v_cnt >= bagel1_y+20 && v_cnt <= bagel1_y+24)||(h_cnt >= bagel1_x+6 && h_cnt <= bagel1_x+8 && v_cnt >= bagel1_y+22 && v_cnt <= bagel1_y+24)||(h_cnt >= bagel1_x+32 && h_cnt <= bagel1_x+34 && v_cnt >= bagel1_y+24 && v_cnt <= bagel1_y+28)||(h_cnt >= bagel1_x+34 && h_cnt <= bagel1_x+36 && v_cnt >= bagel1_y+22 && v_cnt <= bagel1_y+24))
					{vgaRed, vgaGreen, vgaBlue} = 12'hf48; // dark pink
				else if((h_cnt >= bagel1_x+4 && h_cnt <= bagel1_x+6 && v_cnt >= bagel1_y+24 && v_cnt <= bagel1_y+28)||(h_cnt >= bagel1_x+6 && h_cnt <= bagel1_x+8 && v_cnt >= bagel1_y+26 && v_cnt <= bagel1_y+30)||(h_cnt >= bagel1_x+8 && h_cnt <= bagel1_x+12 && v_cnt >= bagel1_y+28 && v_cnt <= bagel1_y+32)||(h_cnt >= bagel1_x+12 && h_cnt <= bagel1_x+26 && v_cnt >= bagel1_y+30 && v_cnt <= bagel1_y+34)||(h_cnt >= bagel1_x+26 && h_cnt <= bagel1_x+30 && v_cnt >= bagel1_y+28 && v_cnt <= bagel1_y+32)||(h_cnt >= bagel1_x+30 && h_cnt <= bagel1_x+32 && v_cnt >= bagel1_y+26 && v_cnt <= bagel1_y+30)||(h_cnt >= bagel1_x+4 && h_cnt <= bagel1_x+6 && v_cnt >= bagel1_y+24 && v_cnt <= bagel1_y+28)||(h_cnt >= bagel1_x+12 && h_cnt <= bagel1_x+14 && v_cnt >= bagel1_y+22 && v_cnt <= bagel1_y+24))
					{vgaRed, vgaGreen, vgaBlue} = 12'hfd5; // yellow
				
				else if((h_cnt >= bagel2_x+12 && h_cnt <= bagel2_x+26 && v_cnt >= bagel2_y && v_cnt <= bagel2_y+2)||(h_cnt >= bagel2_x+8 && h_cnt <= bagel2_x+12 && v_cnt >= bagel2_y+2 && v_cnt <= bagel2_y+4)||(h_cnt >= bagel2_x+26 && h_cnt <= bagel2_x+30 && v_cnt >= bagel2_y+2 && v_cnt <= bagel2_y+4)||(h_cnt >= bagel2_x+6 && h_cnt <= bagel2_x+8 && v_cnt >= bagel2_y+4 && v_cnt <= bagel2_y+6)||(h_cnt >= bagel2_x+30 && h_cnt <= bagel2_x+32 && v_cnt >= bagel2_y+4 && v_cnt <= bagel2_y+6)||(h_cnt >= bagel2_x+4 && h_cnt <= bagel2_x+6 && v_cnt >= bagel2_y+6 && v_cnt <= bagel2_y+8)||(h_cnt >= bagel2_x+32 && h_cnt <= bagel2_x+34 && v_cnt >= bagel2_y+6 && v_cnt <= bagel2_y+8)||(h_cnt >= bagel2_x+2 && h_cnt <= bagel2_x+4 && v_cnt >= bagel2_y+8 && v_cnt <= bagel2_y+12)||(h_cnt >= bagel2_x+34 && h_cnt <= bagel2_x+36 && v_cnt >= bagel2_y+8 && v_cnt <= bagel2_y+12)||(h_cnt >= bagel2_x && h_cnt <= bagel2_x+2 && v_cnt >= bagel2_y+12 && v_cnt <= bagel2_y+24)||(h_cnt >= bagel2_x+36 && h_cnt <= bagel2_x+38 && v_cnt >= bagel2_y+12 && v_cnt <= bagel2_y+24)||(h_cnt >= bagel2_x+2 && h_cnt <= bagel2_x+4 && v_cnt >= bagel2_y+24 && v_cnt <= bagel2_y+28)||(h_cnt >= bagel2_x+34 && h_cnt <= bagel2_x+36 && v_cnt >= bagel2_y+24 && v_cnt <= bagel2_y+28)||(h_cnt >= bagel2_x+4 && h_cnt <= bagel2_x+6 && v_cnt >= bagel2_y+28 && v_cnt <= bagel2_y+30)||(h_cnt >= bagel2_x+32 && h_cnt <= bagel2_x+34 && v_cnt >= bagel2_y+28 && v_cnt <= bagel2_y+30)||(h_cnt >= bagel2_x+6 && h_cnt <= bagel2_x+8 && v_cnt >= bagel2_y+30 && v_cnt <= bagel2_y+32)||(h_cnt >= bagel2_x+30 && h_cnt <= bagel2_x+32 && v_cnt >= bagel2_y+30 && v_cnt <= bagel2_y+32)||(h_cnt >= bagel2_x+8 && h_cnt <= bagel2_x+12 && v_cnt >= bagel2_y+32 && v_cnt <= bagel2_y+34)||(h_cnt >= bagel2_x+26 && h_cnt <= bagel2_x+30 && v_cnt >= bagel2_y+32 && v_cnt <= bagel2_y+34)||(h_cnt >= bagel2_x+12 && h_cnt <= bagel2_x+26 && v_cnt >= bagel2_y+34 && v_cnt <= bagel2_y+36)||(h_cnt >= bagel2_x+18 && h_cnt <= bagel2_x+22 && v_cnt >= bagel2_y+14 && v_cnt <= bagel2_y+16)||(h_cnt >= bagel2_x+18 && h_cnt <= bagel2_x+22 && v_cnt >= bagel2_y+20 && v_cnt <= bagel2_y+22)||(h_cnt >= bagel2_x+16 && h_cnt <= bagel2_x+18 && v_cnt >= bagel2_y+16 && v_cnt <= bagel2_y+20)||(h_cnt >= bagel2_x+22 && h_cnt <= bagel2_x+24 && v_cnt >= bagel2_y+16 && v_cnt <= bagel2_y+20))
					{vgaRed, vgaGreen, vgaBlue} = 12'h0; // black
				else if((h_cnt >= bagel2_x+14 && h_cnt <= bagel2_x+16 && v_cnt >= bagel2_y+2 && v_cnt <= bagel2_y+4)||(h_cnt >= bagel2_x+24 && h_cnt <= bagel2_x+26 && v_cnt >= bagel2_y+2 && v_cnt <= bagel2_y+4)||(h_cnt >= bagel2_x+8 && h_cnt <= bagel2_x+10 && v_cnt >= bagel2_y+4 && v_cnt <= bagel2_y+6)||(h_cnt >= bagel2_x+26 && h_cnt <= bagel2_x+28 && v_cnt >= bagel2_y+4 && v_cnt <= bagel2_y+6)||(h_cnt >= bagel2_x+6 && h_cnt <= bagel2_x+8 && v_cnt >= bagel2_y+6 && v_cnt <= bagel2_y+8)||(h_cnt >= bagel2_x+14 && h_cnt <= bagel2_x+26 && v_cnt >= bagel2_y+6 && v_cnt <= bagel2_y+8)||(h_cnt >= bagel2_x+28 && h_cnt <= bagel2_x+30 && v_cnt >= bagel2_y+6 && v_cnt <= bagel2_y+8)||(h_cnt >= bagel2_x+4 && h_cnt <= bagel2_x+6 && v_cnt >= bagel2_y+8 && v_cnt <= bagel2_y+10)||(h_cnt >= bagel2_x+12 && h_cnt <= bagel2_x+26 && v_cnt >= bagel2_y+8 && v_cnt <= bagel2_y+10)||(h_cnt >= bagel2_x+28 && h_cnt <= bagel2_x+32 && v_cnt >= bagel2_y+8 && v_cnt <= bagel2_y+10)||(h_cnt >= bagel2_x+10 && h_cnt <= bagel2_x+14 && v_cnt >= bagel2_y+10 && v_cnt <= bagel2_y+20)||(h_cnt >= bagel2_x+24 && h_cnt <= bagel2_x+26 && v_cnt >= bagel2_y+10 && v_cnt <= bagel2_y+14)||(h_cnt >= bagel2_x+30 && h_cnt <= bagel2_x+34 && v_cnt >= bagel2_y+10 && v_cnt <= bagel2_y+18)||(h_cnt >= bagel2_x+28 && h_cnt <= bagel2_x+32 && v_cnt >= bagel2_y+18 && v_cnt <= bagel2_y+20)||(h_cnt >= bagel2_x+4 && h_cnt <= bagel2_x+6 && v_cnt >= bagel2_y+18 && v_cnt <= bagel2_y+20)||(h_cnt >= bagel2_x+6 && h_cnt <= bagel2_x+10 && v_cnt >= bagel2_y+20 && v_cnt <= bagel2_y+22)||(h_cnt >= bagel2_x+12 && h_cnt <= bagel2_x+16 && v_cnt >= bagel2_y+20 && v_cnt <= bagel2_y+22)||(h_cnt >= bagel2_x+26 && h_cnt <= bagel2_x+30 && v_cnt >= bagel2_y+20 && v_cnt <= bagel2_y+22)||(h_cnt >= bagel2_x+34 && h_cnt <= bagel2_x+36 && v_cnt >= bagel2_y+20 && v_cnt <= bagel2_y+22)||(h_cnt >= bagel2_x+4 && h_cnt <= bagel2_x+6 && v_cnt >= bagel2_y+22 && v_cnt <= bagel2_y+24)||(h_cnt >= bagel2_x+8 && h_cnt <= bagel2_x+12 && v_cnt >= bagel2_y+22 && v_cnt <= bagel2_y+24)||(h_cnt >= bagel2_x+14 && h_cnt <= bagel2_x+22 && v_cnt >= bagel2_y+22 && v_cnt <= bagel2_y+24)||(h_cnt >= bagel2_x+24 && h_cnt <= bagel2_x+28 && v_cnt >= bagel2_y+22 && v_cnt <= bagel2_y+24)||(h_cnt >= bagel2_x+32 && h_cnt <= bagel2_x+34 && v_cnt >= bagel2_y+22 && v_cnt <= bagel2_y+24)||(h_cnt >= bagel2_x+6 && h_cnt <= bagel2_x+8 && v_cnt >= bagel2_y+24 && v_cnt <= bagel2_y+26)||(h_cnt >= bagel2_x+12 && h_cnt <= bagel2_x+24 && v_cnt >= bagel2_y+24 && v_cnt <= bagel2_y+26)||(h_cnt >= bagel2_x+30 && h_cnt <= bagel2_x+32 && v_cnt >= bagel2_y+24 && v_cnt <= bagel2_y+26)||(h_cnt >= bagel2_x+8 && h_cnt <= bagel2_x+10 && v_cnt >= bagel2_y+26 && v_cnt <= bagel2_y+28)||(h_cnt >= bagel2_x+28 && h_cnt <= bagel2_x+30 && v_cnt >= bagel2_y+26 && v_cnt <= bagel2_y+28)||(h_cnt >= bagel2_x+12 && h_cnt <= bagel2_x+14 && v_cnt >= bagel2_y+28 && v_cnt <= bagel2_y+30)||(h_cnt >= bagel2_x+24 && h_cnt <= bagel2_x+26 && v_cnt >= bagel2_y+28 && v_cnt <= bagel2_y+30))
					{vgaRed, vgaGreen, vgaBlue} = 12'hf9c; // baby pink
				else if((h_cnt >= bagel2_x+16 && h_cnt <= bagel2_x+24 && v_cnt >= bagel2_y+2 && v_cnt <= bagel2_y+4)||(h_cnt >= bagel2_x+10 && h_cnt <= bagel2_x+26 && v_cnt >= bagel2_y+4 && v_cnt <= bagel2_y+6)||(h_cnt >= bagel2_x+8 && h_cnt <= bagel2_x+14 && v_cnt >= bagel2_y+6 && v_cnt <= bagel2_y+8)||(h_cnt >= bagel2_x+26 && h_cnt <= bagel2_x+28 && v_cnt >= bagel2_y+6 && v_cnt <= bagel2_y+20)||(h_cnt >= bagel2_x+28 && h_cnt <= bagel2_x+30 && v_cnt >= bagel2_y+10 && v_cnt <= bagel2_y+18)||(h_cnt >= bagel2_x+24 && h_cnt <= bagel2_x+26 && v_cnt >= bagel2_y+14 && v_cnt <= bagel2_y+22)||(h_cnt >= bagel2_x+14 && h_cnt <= bagel2_x+24 && v_cnt >= bagel2_y+10 && v_cnt <= bagel2_y+14)||(h_cnt >= bagel2_x+4 && h_cnt <= bagel2_x+10 && v_cnt >= bagel2_y+10 && v_cnt <= bagel2_y+18)||(h_cnt >= bagel2_x+2 && h_cnt <= bagel2_x+4 && v_cnt >= bagel2_y+12 && v_cnt <= bagel2_y+24)||(h_cnt >= bagel2_x+6 && h_cnt <= bagel2_x+10 && v_cnt >= bagel2_y+18 && v_cnt <= bagel2_y+20)||(h_cnt >= bagel2_x+4 && h_cnt <= bagel2_x+6 && v_cnt >= bagel2_y+20 && v_cnt <= bagel2_y+22)||(h_cnt >= bagel2_x+34 && h_cnt <= bagel2_x+36 && v_cnt >= bagel2_y+12 && v_cnt <= bagel2_y+20)||(h_cnt >= bagel2_x+22 && h_cnt <= bagel2_x+24 && v_cnt >= bagel2_y+14 && v_cnt <= bagel2_y+16)||(h_cnt >= bagel2_x+14 && h_cnt <= bagel2_x+18 && v_cnt >= bagel2_y+14 && v_cnt <= bagel2_y+16)||(h_cnt >= bagel2_x+14 && h_cnt <= bagel2_x+16 && v_cnt >= bagel2_y+16 && v_cnt <= bagel2_y+20)||(h_cnt >= bagel2_x+32 && h_cnt <= bagel2_x+34 && v_cnt >= bagel2_y+18 && v_cnt <= bagel2_y+22)||(h_cnt >= bagel2_x+30 && h_cnt <= bagel2_x+32 && v_cnt >= bagel2_y+20 && v_cnt <= bagel2_y+24)||(h_cnt >= bagel2_x+28 && h_cnt <= bagel2_x+30 && v_cnt >= bagel2_y+22 && v_cnt <= bagel2_y+26)||(h_cnt >= bagel2_x+24 && h_cnt <= bagel2_x+28 && v_cnt >= bagel2_y+24 && v_cnt <= bagel2_y+28)||(h_cnt >= bagel2_x+14 && h_cnt <= bagel2_x+26 && v_cnt >= bagel2_y+26 && v_cnt <= bagel2_y+30)||(h_cnt >= bagel2_x+10 && h_cnt <= bagel2_x+14 && v_cnt >= bagel2_y+26 && v_cnt <= bagel2_y+28)||(h_cnt >= bagel2_x+8 && h_cnt <= bagel2_x+12 && v_cnt >= bagel2_y+24 && v_cnt <= bagel2_y+26)||(h_cnt >= bagel2_x+6 && h_cnt <= bagel2_x+12 && v_cnt >= bagel2_y+8 && v_cnt <= bagel2_y+10))
					{vgaRed, vgaGreen, vgaBlue} = 12'hf69; // light pink
				else if((h_cnt >= bagel2_x+12 && h_cnt <= bagel2_x+14 && v_cnt >= bagel2_y+2 && v_cnt <= bagel2_y+4)||(h_cnt >= bagel2_x+28 && h_cnt <= bagel2_x+30 && v_cnt >= bagel2_y+4 && v_cnt <= bagel2_y+6)||(h_cnt >= bagel2_x+30 && h_cnt <= bagel2_x+32 && v_cnt >= bagel2_y+6 && v_cnt <= bagel2_y+8)||(h_cnt >= bagel2_x+32 && h_cnt <= bagel2_x+34 && v_cnt >= bagel2_y+8 && v_cnt <= bagel2_y+10)||(h_cnt >= bagel2_x+10 && h_cnt <= bagel2_x+12 && v_cnt >= bagel2_y+20 && v_cnt <= bagel2_y+22)||(h_cnt >= bagel2_x+16 && h_cnt <= bagel2_x+18 && v_cnt >= bagel2_y+20 && v_cnt <= bagel2_y+22)||(h_cnt >= bagel2_x+22 && h_cnt <= bagel2_x+24 && v_cnt >= bagel2_y+20 && v_cnt <= bagel2_y+24)||(h_cnt >= bagel2_x+6 && h_cnt <= bagel2_x+8 && v_cnt >= bagel2_y+22 && v_cnt <= bagel2_y+24)||(h_cnt >= bagel2_x+32 && h_cnt <= bagel2_x+34 && v_cnt >= bagel2_y+24 && v_cnt <= bagel2_y+28)||(h_cnt >= bagel2_x+34 && h_cnt <= bagel2_x+36 && v_cnt >= bagel2_y+22 && v_cnt <= bagel2_y+24))
					{vgaRed, vgaGreen, vgaBlue} = 12'hf48; // dark pink
				else if((h_cnt >= bagel2_x+4 && h_cnt <= bagel2_x+6 && v_cnt >= bagel2_y+24 && v_cnt <= bagel2_y+28)||(h_cnt >= bagel2_x+6 && h_cnt <= bagel2_x+8 && v_cnt >= bagel2_y+26 && v_cnt <= bagel2_y+30)||(h_cnt >= bagel2_x+8 && h_cnt <= bagel2_x+12 && v_cnt >= bagel2_y+28 && v_cnt <= bagel2_y+32)||(h_cnt >= bagel2_x+12 && h_cnt <= bagel2_x+26 && v_cnt >= bagel2_y+30 && v_cnt <= bagel2_y+34)||(h_cnt >= bagel2_x+26 && h_cnt <= bagel2_x+30 && v_cnt >= bagel2_y+28 && v_cnt <= bagel2_y+32)||(h_cnt >= bagel2_x+30 && h_cnt <= bagel2_x+32 && v_cnt >= bagel2_y+26 && v_cnt <= bagel2_y+30)||(h_cnt >= bagel2_x+4 && h_cnt <= bagel2_x+6 && v_cnt >= bagel2_y+24 && v_cnt <= bagel2_y+28)||(h_cnt >= bagel2_x+12 && h_cnt <= bagel2_x+14 && v_cnt >= bagel2_y+22 && v_cnt <= bagel2_y+24))
					{vgaRed, vgaGreen, vgaBlue} = 12'hfd5; // yellow
				
				else if((h_cnt >= bagel3_x+12 && h_cnt <= bagel3_x+26 && v_cnt >= bagel3_y && v_cnt <= bagel3_y+2)||(h_cnt >= bagel3_x+8 && h_cnt <= bagel3_x+12 && v_cnt >= bagel3_y+2 && v_cnt <= bagel3_y+4)||(h_cnt >= bagel3_x+26 && h_cnt <= bagel3_x+30 && v_cnt >= bagel3_y+2 && v_cnt <= bagel3_y+4)||(h_cnt >= bagel3_x+6 && h_cnt <= bagel3_x+8 && v_cnt >= bagel3_y+4 && v_cnt <= bagel3_y+6)||(h_cnt >= bagel3_x+30 && h_cnt <= bagel3_x+32 && v_cnt >= bagel3_y+4 && v_cnt <= bagel3_y+6)||(h_cnt >= bagel3_x+4 && h_cnt <= bagel3_x+6 && v_cnt >= bagel3_y+6 && v_cnt <= bagel3_y+8)||(h_cnt >= bagel3_x+32 && h_cnt <= bagel3_x+34 && v_cnt >= bagel3_y+6 && v_cnt <= bagel3_y+8)||(h_cnt >= bagel3_x+2 && h_cnt <= bagel3_x+4 && v_cnt >= bagel3_y+8 && v_cnt <= bagel3_y+12)||(h_cnt >= bagel3_x+34 && h_cnt <= bagel3_x+36 && v_cnt >= bagel3_y+8 && v_cnt <= bagel3_y+12)||(h_cnt >= bagel3_x && h_cnt <= bagel3_x+2 && v_cnt >= bagel3_y+12 && v_cnt <= bagel3_y+24)||(h_cnt >= bagel3_x+36 && h_cnt <= bagel3_x+38 && v_cnt >= bagel3_y+12 && v_cnt <= bagel3_y+24)||(h_cnt >= bagel3_x+2 && h_cnt <= bagel3_x+4 && v_cnt >= bagel3_y+24 && v_cnt <= bagel3_y+28)||(h_cnt >= bagel3_x+34 && h_cnt <= bagel3_x+36 && v_cnt >= bagel3_y+24 && v_cnt <= bagel3_y+28)||(h_cnt >= bagel3_x+4 && h_cnt <= bagel3_x+6 && v_cnt >= bagel3_y+28 && v_cnt <= bagel3_y+30)||(h_cnt >= bagel3_x+32 && h_cnt <= bagel3_x+34 && v_cnt >= bagel3_y+28 && v_cnt <= bagel3_y+30)||(h_cnt >= bagel3_x+6 && h_cnt <= bagel3_x+8 && v_cnt >= bagel3_y+30 && v_cnt <= bagel3_y+32)||(h_cnt >= bagel3_x+30 && h_cnt <= bagel3_x+32 && v_cnt >= bagel3_y+30 && v_cnt <= bagel3_y+32)||(h_cnt >= bagel3_x+8 && h_cnt <= bagel3_x+12 && v_cnt >= bagel3_y+32 && v_cnt <= bagel3_y+34)||(h_cnt >= bagel3_x+26 && h_cnt <= bagel3_x+30 && v_cnt >= bagel3_y+32 && v_cnt <= bagel3_y+34)||(h_cnt >= bagel3_x+12 && h_cnt <= bagel3_x+26 && v_cnt >= bagel3_y+34 && v_cnt <= bagel3_y+36)||(h_cnt >= bagel3_x+18 && h_cnt <= bagel3_x+22 && v_cnt >= bagel3_y+14 && v_cnt <= bagel3_y+16)||(h_cnt >= bagel3_x+18 && h_cnt <= bagel3_x+22 && v_cnt >= bagel3_y+20 && v_cnt <= bagel3_y+22)||(h_cnt >= bagel3_x+16 && h_cnt <= bagel3_x+18 && v_cnt >= bagel3_y+16 && v_cnt <= bagel3_y+20)||(h_cnt >= bagel3_x+22 && h_cnt <= bagel3_x+24 && v_cnt >= bagel3_y+16 && v_cnt <= bagel3_y+20))
					{vgaRed, vgaGreen, vgaBlue} = 12'h0; // black
				else if((h_cnt >= bagel3_x+14 && h_cnt <= bagel3_x+16 && v_cnt >= bagel3_y+2 && v_cnt <= bagel3_y+4)||(h_cnt >= bagel3_x+24 && h_cnt <= bagel3_x+26 && v_cnt >= bagel3_y+2 && v_cnt <= bagel3_y+4)||(h_cnt >= bagel3_x+8 && h_cnt <= bagel3_x+10 && v_cnt >= bagel3_y+4 && v_cnt <= bagel3_y+6)||(h_cnt >= bagel3_x+26 && h_cnt <= bagel3_x+28 && v_cnt >= bagel3_y+4 && v_cnt <= bagel3_y+6)||(h_cnt >= bagel3_x+6 && h_cnt <= bagel3_x+8 && v_cnt >= bagel3_y+6 && v_cnt <= bagel3_y+8)||(h_cnt >= bagel3_x+14 && h_cnt <= bagel3_x+26 && v_cnt >= bagel3_y+6 && v_cnt <= bagel3_y+8)||(h_cnt >= bagel3_x+28 && h_cnt <= bagel3_x+30 && v_cnt >= bagel3_y+6 && v_cnt <= bagel3_y+8)||(h_cnt >= bagel3_x+4 && h_cnt <= bagel3_x+6 && v_cnt >= bagel3_y+8 && v_cnt <= bagel3_y+10)||(h_cnt >= bagel3_x+12 && h_cnt <= bagel3_x+26 && v_cnt >= bagel3_y+8 && v_cnt <= bagel3_y+10)||(h_cnt >= bagel3_x+28 && h_cnt <= bagel3_x+32 && v_cnt >= bagel3_y+8 && v_cnt <= bagel3_y+10)||(h_cnt >= bagel3_x+10 && h_cnt <= bagel3_x+14 && v_cnt >= bagel3_y+10 && v_cnt <= bagel3_y+20)||(h_cnt >= bagel3_x+24 && h_cnt <= bagel3_x+26 && v_cnt >= bagel3_y+10 && v_cnt <= bagel3_y+14)||(h_cnt >= bagel3_x+30 && h_cnt <= bagel3_x+34 && v_cnt >= bagel3_y+10 && v_cnt <= bagel3_y+18)||(h_cnt >= bagel3_x+28 && h_cnt <= bagel3_x+32 && v_cnt >= bagel3_y+18 && v_cnt <= bagel3_y+20)||(h_cnt >= bagel3_x+4 && h_cnt <= bagel3_x+6 && v_cnt >= bagel3_y+18 && v_cnt <= bagel3_y+20)||(h_cnt >= bagel3_x+6 && h_cnt <= bagel3_x+10 && v_cnt >= bagel3_y+20 && v_cnt <= bagel3_y+22)||(h_cnt >= bagel3_x+12 && h_cnt <= bagel3_x+16 && v_cnt >= bagel3_y+20 && v_cnt <= bagel3_y+22)||(h_cnt >= bagel3_x+26 && h_cnt <= bagel3_x+30 && v_cnt >= bagel3_y+20 && v_cnt <= bagel3_y+22)||(h_cnt >= bagel3_x+34 && h_cnt <= bagel3_x+36 && v_cnt >= bagel3_y+20 && v_cnt <= bagel3_y+22)||(h_cnt >= bagel3_x+4 && h_cnt <= bagel3_x+6 && v_cnt >= bagel3_y+22 && v_cnt <= bagel3_y+24)||(h_cnt >= bagel3_x+8 && h_cnt <= bagel3_x+12 && v_cnt >= bagel3_y+22 && v_cnt <= bagel3_y+24)||(h_cnt >= bagel3_x+14 && h_cnt <= bagel3_x+22 && v_cnt >= bagel3_y+22 && v_cnt <= bagel3_y+24)||(h_cnt >= bagel3_x+24 && h_cnt <= bagel3_x+28 && v_cnt >= bagel3_y+22 && v_cnt <= bagel3_y+24)||(h_cnt >= bagel3_x+32 && h_cnt <= bagel3_x+34 && v_cnt >= bagel3_y+22 && v_cnt <= bagel3_y+24)||(h_cnt >= bagel3_x+6 && h_cnt <= bagel3_x+8 && v_cnt >= bagel3_y+24 && v_cnt <= bagel3_y+26)||(h_cnt >= bagel3_x+12 && h_cnt <= bagel3_x+24 && v_cnt >= bagel3_y+24 && v_cnt <= bagel3_y+26)||(h_cnt >= bagel3_x+30 && h_cnt <= bagel3_x+32 && v_cnt >= bagel3_y+24 && v_cnt <= bagel3_y+26)||(h_cnt >= bagel3_x+8 && h_cnt <= bagel3_x+10 && v_cnt >= bagel3_y+26 && v_cnt <= bagel3_y+28)||(h_cnt >= bagel3_x+28 && h_cnt <= bagel3_x+30 && v_cnt >= bagel3_y+26 && v_cnt <= bagel3_y+28)||(h_cnt >= bagel3_x+12 && h_cnt <= bagel3_x+14 && v_cnt >= bagel3_y+28 && v_cnt <= bagel3_y+30)||(h_cnt >= bagel3_x+24 && h_cnt <= bagel3_x+26 && v_cnt >= bagel3_y+28 && v_cnt <= bagel3_y+30))
					{vgaRed, vgaGreen, vgaBlue} = 12'hf9c; // baby pink
				else if((h_cnt >= bagel3_x+16 && h_cnt <= bagel3_x+24 && v_cnt >= bagel3_y+2 && v_cnt <= bagel3_y+4)||(h_cnt >= bagel3_x+10 && h_cnt <= bagel3_x+26 && v_cnt >= bagel3_y+4 && v_cnt <= bagel3_y+6)||(h_cnt >= bagel3_x+8 && h_cnt <= bagel3_x+14 && v_cnt >= bagel3_y+6 && v_cnt <= bagel3_y+8)||(h_cnt >= bagel3_x+26 && h_cnt <= bagel3_x+28 && v_cnt >= bagel3_y+6 && v_cnt <= bagel3_y+20)||(h_cnt >= bagel3_x+28 && h_cnt <= bagel3_x+30 && v_cnt >= bagel3_y+10 && v_cnt <= bagel3_y+18)||(h_cnt >= bagel3_x+24 && h_cnt <= bagel3_x+26 && v_cnt >= bagel3_y+14 && v_cnt <= bagel3_y+22)||(h_cnt >= bagel3_x+14 && h_cnt <= bagel3_x+24 && v_cnt >= bagel3_y+10 && v_cnt <= bagel3_y+14)||(h_cnt >= bagel3_x+4 && h_cnt <= bagel3_x+10 && v_cnt >= bagel3_y+10 && v_cnt <= bagel3_y+18)||(h_cnt >= bagel3_x+2 && h_cnt <= bagel3_x+4 && v_cnt >= bagel3_y+12 && v_cnt <= bagel3_y+24)||(h_cnt >= bagel3_x+6 && h_cnt <= bagel3_x+10 && v_cnt >= bagel3_y+18 && v_cnt <= bagel3_y+20)||(h_cnt >= bagel3_x+4 && h_cnt <= bagel3_x+6 && v_cnt >= bagel3_y+20 && v_cnt <= bagel3_y+22)||(h_cnt >= bagel3_x+34 && h_cnt <= bagel3_x+36 && v_cnt >= bagel3_y+12 && v_cnt <= bagel3_y+20)||(h_cnt >= bagel3_x+22 && h_cnt <= bagel3_x+24 && v_cnt >= bagel3_y+14 && v_cnt <= bagel3_y+16)||(h_cnt >= bagel3_x+14 && h_cnt <= bagel3_x+18 && v_cnt >= bagel3_y+14 && v_cnt <= bagel3_y+16)||(h_cnt >= bagel3_x+14 && h_cnt <= bagel3_x+16 && v_cnt >= bagel3_y+16 && v_cnt <= bagel3_y+20)||(h_cnt >= bagel3_x+32 && h_cnt <= bagel3_x+34 && v_cnt >= bagel3_y+18 && v_cnt <= bagel3_y+22)||(h_cnt >= bagel3_x+30 && h_cnt <= bagel3_x+32 && v_cnt >= bagel3_y+20 && v_cnt <= bagel3_y+24)||(h_cnt >= bagel3_x+28 && h_cnt <= bagel3_x+30 && v_cnt >= bagel3_y+22 && v_cnt <= bagel3_y+26)||(h_cnt >= bagel3_x+24 && h_cnt <= bagel3_x+28 && v_cnt >= bagel3_y+24 && v_cnt <= bagel3_y+28)||(h_cnt >= bagel3_x+14 && h_cnt <= bagel3_x+26 && v_cnt >= bagel3_y+26 && v_cnt <= bagel3_y+30)||(h_cnt >= bagel3_x+10 && h_cnt <= bagel3_x+14 && v_cnt >= bagel3_y+26 && v_cnt <= bagel3_y+28)||(h_cnt >= bagel3_x+8 && h_cnt <= bagel3_x+12 && v_cnt >= bagel3_y+24 && v_cnt <= bagel3_y+26)||(h_cnt >= bagel3_x+6 && h_cnt <= bagel3_x+12 && v_cnt >= bagel3_y+8 && v_cnt <= bagel3_y+10))
					{vgaRed, vgaGreen, vgaBlue} = 12'hf69; // light pink
				else if((h_cnt >= bagel3_x+12 && h_cnt <= bagel3_x+14 && v_cnt >= bagel3_y+2 && v_cnt <= bagel3_y+4)||(h_cnt >= bagel3_x+28 && h_cnt <= bagel3_x+30 && v_cnt >= bagel3_y+4 && v_cnt <= bagel3_y+6)||(h_cnt >= bagel3_x+30 && h_cnt <= bagel3_x+32 && v_cnt >= bagel3_y+6 && v_cnt <= bagel3_y+8)||(h_cnt >= bagel3_x+32 && h_cnt <= bagel3_x+34 && v_cnt >= bagel3_y+8 && v_cnt <= bagel3_y+10)||(h_cnt >= bagel3_x+10 && h_cnt <= bagel3_x+12 && v_cnt >= bagel3_y+20 && v_cnt <= bagel3_y+22)||(h_cnt >= bagel3_x+16 && h_cnt <= bagel3_x+18 && v_cnt >= bagel3_y+20 && v_cnt <= bagel3_y+22)||(h_cnt >= bagel3_x+22 && h_cnt <= bagel3_x+24 && v_cnt >= bagel3_y+20 && v_cnt <= bagel3_y+24)||(h_cnt >= bagel3_x+6 && h_cnt <= bagel3_x+8 && v_cnt >= bagel3_y+22 && v_cnt <= bagel3_y+24)||(h_cnt >= bagel3_x+32 && h_cnt <= bagel3_x+34 && v_cnt >= bagel3_y+24 && v_cnt <= bagel3_y+28)||(h_cnt >= bagel3_x+34 && h_cnt <= bagel3_x+36 && v_cnt >= bagel3_y+22 && v_cnt <= bagel3_y+24))
					{vgaRed, vgaGreen, vgaBlue} = 12'hf48; // dark pink
				else if((h_cnt >= bagel3_x+4 && h_cnt <= bagel3_x+6 && v_cnt >= bagel3_y+24 && v_cnt <= bagel3_y+28)||(h_cnt >= bagel3_x+6 && h_cnt <= bagel3_x+8 && v_cnt >= bagel3_y+26 && v_cnt <= bagel3_y+30)||(h_cnt >= bagel3_x+8 && h_cnt <= bagel3_x+12 && v_cnt >= bagel3_y+28 && v_cnt <= bagel3_y+32)||(h_cnt >= bagel3_x+12 && h_cnt <= bagel3_x+26 && v_cnt >= bagel3_y+30 && v_cnt <= bagel3_y+34)||(h_cnt >= bagel3_x+26 && h_cnt <= bagel3_x+30 && v_cnt >= bagel3_y+28 && v_cnt <= bagel3_y+32)||(h_cnt >= bagel3_x+30 && h_cnt <= bagel3_x+32 && v_cnt >= bagel3_y+26 && v_cnt <= bagel3_y+30)||(h_cnt >= bagel3_x+4 && h_cnt <= bagel3_x+6 && v_cnt >= bagel3_y+24 && v_cnt <= bagel3_y+28)||(h_cnt >= bagel3_x+12 && h_cnt <= bagel3_x+14 && v_cnt >= bagel3_y+22 && v_cnt <= bagel3_y+24))
					{vgaRed, vgaGreen, vgaBlue} = 12'hfd5; // yellow
				
				else if((h_cnt >= bagel4_x+12 && h_cnt <= bagel4_x+26 && v_cnt >= bagel4_y && v_cnt <= bagel4_y+2)||(h_cnt >= bagel4_x+8 && h_cnt <= bagel4_x+12 && v_cnt >= bagel4_y+2 && v_cnt <= bagel4_y+4)||(h_cnt >= bagel4_x+26 && h_cnt <= bagel4_x+30 && v_cnt >= bagel4_y+2 && v_cnt <= bagel4_y+4)||(h_cnt >= bagel4_x+6 && h_cnt <= bagel4_x+8 && v_cnt >= bagel4_y+4 && v_cnt <= bagel4_y+6)||(h_cnt >= bagel4_x+30 && h_cnt <= bagel4_x+32 && v_cnt >= bagel4_y+4 && v_cnt <= bagel4_y+6)||(h_cnt >= bagel4_x+4 && h_cnt <= bagel4_x+6 && v_cnt >= bagel4_y+6 && v_cnt <= bagel4_y+8)||(h_cnt >= bagel4_x+32 && h_cnt <= bagel4_x+34 && v_cnt >= bagel4_y+6 && v_cnt <= bagel4_y+8)||(h_cnt >= bagel4_x+2 && h_cnt <= bagel4_x+4 && v_cnt >= bagel4_y+8 && v_cnt <= bagel4_y+12)||(h_cnt >= bagel4_x+34 && h_cnt <= bagel4_x+36 && v_cnt >= bagel4_y+8 && v_cnt <= bagel4_y+12)||(h_cnt >= bagel4_x && h_cnt <= bagel4_x+2 && v_cnt >= bagel4_y+12 && v_cnt <= bagel4_y+24)||(h_cnt >= bagel4_x+36 && h_cnt <= bagel4_x+38 && v_cnt >= bagel4_y+12 && v_cnt <= bagel4_y+24)||(h_cnt >= bagel4_x+2 && h_cnt <= bagel4_x+4 && v_cnt >= bagel4_y+24 && v_cnt <= bagel4_y+28)||(h_cnt >= bagel4_x+34 && h_cnt <= bagel4_x+36 && v_cnt >= bagel4_y+24 && v_cnt <= bagel4_y+28)||(h_cnt >= bagel4_x+4 && h_cnt <= bagel4_x+6 && v_cnt >= bagel4_y+28 && v_cnt <= bagel4_y+30)||(h_cnt >= bagel4_x+32 && h_cnt <= bagel4_x+34 && v_cnt >= bagel4_y+28 && v_cnt <= bagel4_y+30)||(h_cnt >= bagel4_x+6 && h_cnt <= bagel4_x+8 && v_cnt >= bagel4_y+30 && v_cnt <= bagel4_y+32)||(h_cnt >= bagel4_x+30 && h_cnt <= bagel4_x+32 && v_cnt >= bagel4_y+30 && v_cnt <= bagel4_y+32)||(h_cnt >= bagel4_x+8 && h_cnt <= bagel4_x+12 && v_cnt >= bagel4_y+32 && v_cnt <= bagel4_y+34)||(h_cnt >= bagel4_x+26 && h_cnt <= bagel4_x+30 && v_cnt >= bagel4_y+32 && v_cnt <= bagel4_y+34)||(h_cnt >= bagel4_x+12 && h_cnt <= bagel4_x+26 && v_cnt >= bagel4_y+34 && v_cnt <= bagel4_y+36)||(h_cnt >= bagel4_x+18 && h_cnt <= bagel4_x+22 && v_cnt >= bagel4_y+14 && v_cnt <= bagel4_y+16)||(h_cnt >= bagel4_x+18 && h_cnt <= bagel4_x+22 && v_cnt >= bagel4_y+20 && v_cnt <= bagel4_y+22)||(h_cnt >= bagel4_x+16 && h_cnt <= bagel4_x+18 && v_cnt >= bagel4_y+16 && v_cnt <= bagel4_y+20)||(h_cnt >= bagel4_x+22 && h_cnt <= bagel4_x+24 && v_cnt >= bagel4_y+16 && v_cnt <= bagel4_y+20))
					{vgaRed, vgaGreen, vgaBlue} = 12'h0; // black
				else if((h_cnt >= bagel4_x+14 && h_cnt <= bagel4_x+16 && v_cnt >= bagel4_y+2 && v_cnt <= bagel4_y+4)||(h_cnt >= bagel4_x+24 && h_cnt <= bagel4_x+26 && v_cnt >= bagel4_y+2 && v_cnt <= bagel4_y+4)||(h_cnt >= bagel4_x+8 && h_cnt <= bagel4_x+10 && v_cnt >= bagel4_y+4 && v_cnt <= bagel4_y+6)||(h_cnt >= bagel4_x+26 && h_cnt <= bagel4_x+28 && v_cnt >= bagel4_y+4 && v_cnt <= bagel4_y+6)||(h_cnt >= bagel4_x+6 && h_cnt <= bagel4_x+8 && v_cnt >= bagel4_y+6 && v_cnt <= bagel4_y+8)||(h_cnt >= bagel4_x+14 && h_cnt <= bagel4_x+26 && v_cnt >= bagel4_y+6 && v_cnt <= bagel4_y+8)||(h_cnt >= bagel4_x+28 && h_cnt <= bagel4_x+30 && v_cnt >= bagel4_y+6 && v_cnt <= bagel4_y+8)||(h_cnt >= bagel4_x+4 && h_cnt <= bagel4_x+6 && v_cnt >= bagel4_y+8 && v_cnt <= bagel4_y+10)||(h_cnt >= bagel4_x+12 && h_cnt <= bagel4_x+26 && v_cnt >= bagel4_y+8 && v_cnt <= bagel4_y+10)||(h_cnt >= bagel4_x+28 && h_cnt <= bagel4_x+32 && v_cnt >= bagel4_y+8 && v_cnt <= bagel4_y+10)||(h_cnt >= bagel4_x+10 && h_cnt <= bagel4_x+14 && v_cnt >= bagel4_y+10 && v_cnt <= bagel4_y+20)||(h_cnt >= bagel4_x+24 && h_cnt <= bagel4_x+26 && v_cnt >= bagel4_y+10 && v_cnt <= bagel4_y+14)||(h_cnt >= bagel4_x+30 && h_cnt <= bagel4_x+34 && v_cnt >= bagel4_y+10 && v_cnt <= bagel4_y+18)||(h_cnt >= bagel4_x+28 && h_cnt <= bagel4_x+32 && v_cnt >= bagel4_y+18 && v_cnt <= bagel4_y+20)||(h_cnt >= bagel4_x+4 && h_cnt <= bagel4_x+6 && v_cnt >= bagel4_y+18 && v_cnt <= bagel4_y+20)||(h_cnt >= bagel4_x+6 && h_cnt <= bagel4_x+10 && v_cnt >= bagel4_y+20 && v_cnt <= bagel4_y+22)||(h_cnt >= bagel4_x+12 && h_cnt <= bagel4_x+16 && v_cnt >= bagel4_y+20 && v_cnt <= bagel4_y+22)||(h_cnt >= bagel4_x+26 && h_cnt <= bagel4_x+30 && v_cnt >= bagel4_y+20 && v_cnt <= bagel4_y+22)||(h_cnt >= bagel4_x+34 && h_cnt <= bagel4_x+36 && v_cnt >= bagel4_y+20 && v_cnt <= bagel4_y+22)||(h_cnt >= bagel4_x+4 && h_cnt <= bagel4_x+6 && v_cnt >= bagel4_y+22 && v_cnt <= bagel4_y+24)||(h_cnt >= bagel4_x+8 && h_cnt <= bagel4_x+12 && v_cnt >= bagel4_y+22 && v_cnt <= bagel4_y+24)||(h_cnt >= bagel4_x+14 && h_cnt <= bagel4_x+22 && v_cnt >= bagel4_y+22 && v_cnt <= bagel4_y+24)||(h_cnt >= bagel4_x+24 && h_cnt <= bagel4_x+28 && v_cnt >= bagel4_y+22 && v_cnt <= bagel4_y+24)||(h_cnt >= bagel4_x+32 && h_cnt <= bagel4_x+34 && v_cnt >= bagel4_y+22 && v_cnt <= bagel4_y+24)||(h_cnt >= bagel4_x+6 && h_cnt <= bagel4_x+8 && v_cnt >= bagel4_y+24 && v_cnt <= bagel4_y+26)||(h_cnt >= bagel4_x+12 && h_cnt <= bagel4_x+24 && v_cnt >= bagel4_y+24 && v_cnt <= bagel4_y+26)||(h_cnt >= bagel4_x+30 && h_cnt <= bagel4_x+32 && v_cnt >= bagel4_y+24 && v_cnt <= bagel4_y+26)||(h_cnt >= bagel4_x+8 && h_cnt <= bagel4_x+10 && v_cnt >= bagel4_y+26 && v_cnt <= bagel4_y+28)||(h_cnt >= bagel4_x+28 && h_cnt <= bagel4_x+30 && v_cnt >= bagel4_y+26 && v_cnt <= bagel4_y+28)||(h_cnt >= bagel4_x+12 && h_cnt <= bagel4_x+14 && v_cnt >= bagel4_y+28 && v_cnt <= bagel4_y+30)||(h_cnt >= bagel4_x+24 && h_cnt <= bagel4_x+26 && v_cnt >= bagel4_y+28 && v_cnt <= bagel4_y+30))
					{vgaRed, vgaGreen, vgaBlue} = 12'hf9c; // baby pink
				else if((h_cnt >= bagel4_x+16 && h_cnt <= bagel4_x+24 && v_cnt >= bagel4_y+2 && v_cnt <= bagel4_y+4)||(h_cnt >= bagel4_x+10 && h_cnt <= bagel4_x+26 && v_cnt >= bagel4_y+4 && v_cnt <= bagel4_y+6)||(h_cnt >= bagel4_x+8 && h_cnt <= bagel4_x+14 && v_cnt >= bagel4_y+6 && v_cnt <= bagel4_y+8)||(h_cnt >= bagel4_x+26 && h_cnt <= bagel4_x+28 && v_cnt >= bagel4_y+6 && v_cnt <= bagel4_y+20)||(h_cnt >= bagel4_x+28 && h_cnt <= bagel4_x+30 && v_cnt >= bagel4_y+10 && v_cnt <= bagel4_y+18)||(h_cnt >= bagel4_x+24 && h_cnt <= bagel4_x+26 && v_cnt >= bagel4_y+14 && v_cnt <= bagel4_y+22)||(h_cnt >= bagel4_x+14 && h_cnt <= bagel4_x+24 && v_cnt >= bagel4_y+10 && v_cnt <= bagel4_y+14)||(h_cnt >= bagel4_x+4 && h_cnt <= bagel4_x+10 && v_cnt >= bagel4_y+10 && v_cnt <= bagel4_y+18)||(h_cnt >= bagel4_x+2 && h_cnt <= bagel4_x+4 && v_cnt >= bagel4_y+12 && v_cnt <= bagel4_y+24)||(h_cnt >= bagel4_x+6 && h_cnt <= bagel4_x+10 && v_cnt >= bagel4_y+18 && v_cnt <= bagel4_y+20)||(h_cnt >= bagel4_x+4 && h_cnt <= bagel4_x+6 && v_cnt >= bagel4_y+20 && v_cnt <= bagel4_y+22)||(h_cnt >= bagel4_x+34 && h_cnt <= bagel4_x+36 && v_cnt >= bagel4_y+12 && v_cnt <= bagel4_y+20)||(h_cnt >= bagel4_x+22 && h_cnt <= bagel4_x+24 && v_cnt >= bagel4_y+14 && v_cnt <= bagel4_y+16)||(h_cnt >= bagel4_x+14 && h_cnt <= bagel4_x+18 && v_cnt >= bagel4_y+14 && v_cnt <= bagel4_y+16)||(h_cnt >= bagel4_x+14 && h_cnt <= bagel4_x+16 && v_cnt >= bagel4_y+16 && v_cnt <= bagel4_y+20)||(h_cnt >= bagel4_x+32 && h_cnt <= bagel4_x+34 && v_cnt >= bagel4_y+18 && v_cnt <= bagel4_y+22)||(h_cnt >= bagel4_x+30 && h_cnt <= bagel4_x+32 && v_cnt >= bagel4_y+20 && v_cnt <= bagel4_y+24)||(h_cnt >= bagel4_x+28 && h_cnt <= bagel4_x+30 && v_cnt >= bagel4_y+22 && v_cnt <= bagel4_y+26)||(h_cnt >= bagel4_x+24 && h_cnt <= bagel4_x+28 && v_cnt >= bagel4_y+24 && v_cnt <= bagel4_y+28)||(h_cnt >= bagel4_x+14 && h_cnt <= bagel4_x+26 && v_cnt >= bagel4_y+26 && v_cnt <= bagel4_y+30)||(h_cnt >= bagel4_x+10 && h_cnt <= bagel4_x+14 && v_cnt >= bagel4_y+26 && v_cnt <= bagel4_y+28)||(h_cnt >= bagel4_x+8 && h_cnt <= bagel4_x+12 && v_cnt >= bagel4_y+24 && v_cnt <= bagel4_y+26)||(h_cnt >= bagel4_x+6 && h_cnt <= bagel4_x+12 && v_cnt >= bagel4_y+8 && v_cnt <= bagel4_y+10))
					{vgaRed, vgaGreen, vgaBlue} = 12'hf69; // light pink
				else if((h_cnt >= bagel4_x+12 && h_cnt <= bagel4_x+14 && v_cnt >= bagel4_y+2 && v_cnt <= bagel4_y+4)||(h_cnt >= bagel4_x+28 && h_cnt <= bagel4_x+30 && v_cnt >= bagel4_y+4 && v_cnt <= bagel4_y+6)||(h_cnt >= bagel4_x+30 && h_cnt <= bagel4_x+32 && v_cnt >= bagel4_y+6 && v_cnt <= bagel4_y+8)||(h_cnt >= bagel4_x+32 && h_cnt <= bagel4_x+34 && v_cnt >= bagel4_y+8 && v_cnt <= bagel4_y+10)||(h_cnt >= bagel4_x+10 && h_cnt <= bagel4_x+12 && v_cnt >= bagel4_y+20 && v_cnt <= bagel4_y+22)||(h_cnt >= bagel4_x+16 && h_cnt <= bagel4_x+18 && v_cnt >= bagel4_y+20 && v_cnt <= bagel4_y+22)||(h_cnt >= bagel4_x+22 && h_cnt <= bagel4_x+24 && v_cnt >= bagel4_y+20 && v_cnt <= bagel4_y+24)||(h_cnt >= bagel4_x+6 && h_cnt <= bagel4_x+8 && v_cnt >= bagel4_y+22 && v_cnt <= bagel4_y+24)||(h_cnt >= bagel4_x+32 && h_cnt <= bagel4_x+34 && v_cnt >= bagel4_y+24 && v_cnt <= bagel4_y+28)||(h_cnt >= bagel4_x+34 && h_cnt <= bagel4_x+36 && v_cnt >= bagel4_y+22 && v_cnt <= bagel4_y+24))
					{vgaRed, vgaGreen, vgaBlue} = 12'hf48; // dark pink
				else if((h_cnt >= bagel4_x+4 && h_cnt <= bagel4_x+6 && v_cnt >= bagel4_y+24 && v_cnt <= bagel4_y+28)||(h_cnt >= bagel4_x+6 && h_cnt <= bagel4_x+8 && v_cnt >= bagel4_y+26 && v_cnt <= bagel4_y+30)||(h_cnt >= bagel4_x+8 && h_cnt <= bagel4_x+12 && v_cnt >= bagel4_y+28 && v_cnt <= bagel4_y+32)||(h_cnt >= bagel4_x+12 && h_cnt <= bagel4_x+26 && v_cnt >= bagel4_y+30 && v_cnt <= bagel4_y+34)||(h_cnt >= bagel4_x+26 && h_cnt <= bagel4_x+30 && v_cnt >= bagel4_y+28 && v_cnt <= bagel4_y+32)||(h_cnt >= bagel4_x+30 && h_cnt <= bagel4_x+32 && v_cnt >= bagel4_y+26 && v_cnt <= bagel4_y+30)||(h_cnt >= bagel4_x+4 && h_cnt <= bagel4_x+6 && v_cnt >= bagel4_y+24 && v_cnt <= bagel4_y+28)||(h_cnt >= bagel4_x+12 && h_cnt <= bagel4_x+14 && v_cnt >= bagel4_y+22 && v_cnt <= bagel4_y+24))
					{vgaRed, vgaGreen, vgaBlue} = 12'hfd5; // yellow
				
				else if((h_cnt >= bagel5_x+12 && h_cnt <= bagel5_x+26 && v_cnt >= bagel5_y && v_cnt <= bagel5_y+2)||(h_cnt >= bagel5_x+8 && h_cnt <= bagel5_x+12 && v_cnt >= bagel5_y+2 && v_cnt <= bagel5_y+4)||(h_cnt >= bagel5_x+26 && h_cnt <= bagel5_x+30 && v_cnt >= bagel5_y+2 && v_cnt <= bagel5_y+4)||(h_cnt >= bagel5_x+6 && h_cnt <= bagel5_x+8 && v_cnt >= bagel5_y+4 && v_cnt <= bagel5_y+6)||(h_cnt >= bagel5_x+30 && h_cnt <= bagel5_x+32 && v_cnt >= bagel5_y+4 && v_cnt <= bagel5_y+6)||(h_cnt >= bagel5_x+4 && h_cnt <= bagel5_x+6 && v_cnt >= bagel5_y+6 && v_cnt <= bagel5_y+8)||(h_cnt >= bagel5_x+32 && h_cnt <= bagel5_x+34 && v_cnt >= bagel5_y+6 && v_cnt <= bagel5_y+8)||(h_cnt >= bagel5_x+2 && h_cnt <= bagel5_x+4 && v_cnt >= bagel5_y+8 && v_cnt <= bagel5_y+12)||(h_cnt >= bagel5_x+34 && h_cnt <= bagel5_x+36 && v_cnt >= bagel5_y+8 && v_cnt <= bagel5_y+12)||(h_cnt >= bagel5_x && h_cnt <= bagel5_x+2 && v_cnt >= bagel5_y+12 && v_cnt <= bagel5_y+24)||(h_cnt >= bagel5_x+36 && h_cnt <= bagel5_x+38 && v_cnt >= bagel5_y+12 && v_cnt <= bagel5_y+24)||(h_cnt >= bagel5_x+2 && h_cnt <= bagel5_x+4 && v_cnt >= bagel5_y+24 && v_cnt <= bagel5_y+28)||(h_cnt >= bagel5_x+34 && h_cnt <= bagel5_x+36 && v_cnt >= bagel5_y+24 && v_cnt <= bagel5_y+28)||(h_cnt >= bagel5_x+4 && h_cnt <= bagel5_x+6 && v_cnt >= bagel5_y+28 && v_cnt <= bagel5_y+30)||(h_cnt >= bagel5_x+32 && h_cnt <= bagel5_x+34 && v_cnt >= bagel5_y+28 && v_cnt <= bagel5_y+30)||(h_cnt >= bagel5_x+6 && h_cnt <= bagel5_x+8 && v_cnt >= bagel5_y+30 && v_cnt <= bagel5_y+32)||(h_cnt >= bagel5_x+30 && h_cnt <= bagel5_x+32 && v_cnt >= bagel5_y+30 && v_cnt <= bagel5_y+32)||(h_cnt >= bagel5_x+8 && h_cnt <= bagel5_x+12 && v_cnt >= bagel5_y+32 && v_cnt <= bagel5_y+34)||(h_cnt >= bagel5_x+26 && h_cnt <= bagel5_x+30 && v_cnt >= bagel5_y+32 && v_cnt <= bagel5_y+34)||(h_cnt >= bagel5_x+12 && h_cnt <= bagel5_x+26 && v_cnt >= bagel5_y+34 && v_cnt <= bagel5_y+36)||(h_cnt >= bagel5_x+18 && h_cnt <= bagel5_x+22 && v_cnt >= bagel5_y+14 && v_cnt <= bagel5_y+16)||(h_cnt >= bagel5_x+18 && h_cnt <= bagel5_x+22 && v_cnt >= bagel5_y+20 && v_cnt <= bagel5_y+22)||(h_cnt >= bagel5_x+16 && h_cnt <= bagel5_x+18 && v_cnt >= bagel5_y+16 && v_cnt <= bagel5_y+20)||(h_cnt >= bagel5_x+22 && h_cnt <= bagel5_x+24 && v_cnt >= bagel5_y+16 && v_cnt <= bagel5_y+20))
					{vgaRed, vgaGreen, vgaBlue} = 12'h0; // black
				else if((h_cnt >= bagel5_x+14 && h_cnt <= bagel5_x+16 && v_cnt >= bagel5_y+2 && v_cnt <= bagel5_y+4)||(h_cnt >= bagel5_x+24 && h_cnt <= bagel5_x+26 && v_cnt >= bagel5_y+2 && v_cnt <= bagel5_y+4)||(h_cnt >= bagel5_x+8 && h_cnt <= bagel5_x+10 && v_cnt >= bagel5_y+4 && v_cnt <= bagel5_y+6)||(h_cnt >= bagel5_x+26 && h_cnt <= bagel5_x+28 && v_cnt >= bagel5_y+4 && v_cnt <= bagel5_y+6)||(h_cnt >= bagel5_x+6 && h_cnt <= bagel5_x+8 && v_cnt >= bagel5_y+6 && v_cnt <= bagel5_y+8)||(h_cnt >= bagel5_x+14 && h_cnt <= bagel5_x+26 && v_cnt >= bagel5_y+6 && v_cnt <= bagel5_y+8)||(h_cnt >= bagel5_x+28 && h_cnt <= bagel5_x+30 && v_cnt >= bagel5_y+6 && v_cnt <= bagel5_y+8)||(h_cnt >= bagel5_x+4 && h_cnt <= bagel5_x+6 && v_cnt >= bagel5_y+8 && v_cnt <= bagel5_y+10)||(h_cnt >= bagel5_x+12 && h_cnt <= bagel5_x+26 && v_cnt >= bagel5_y+8 && v_cnt <= bagel5_y+10)||(h_cnt >= bagel5_x+28 && h_cnt <= bagel5_x+32 && v_cnt >= bagel5_y+8 && v_cnt <= bagel5_y+10)||(h_cnt >= bagel5_x+10 && h_cnt <= bagel5_x+14 && v_cnt >= bagel5_y+10 && v_cnt <= bagel5_y+20)||(h_cnt >= bagel5_x+24 && h_cnt <= bagel5_x+26 && v_cnt >= bagel5_y+10 && v_cnt <= bagel5_y+14)||(h_cnt >= bagel5_x+30 && h_cnt <= bagel5_x+34 && v_cnt >= bagel5_y+10 && v_cnt <= bagel5_y+18)||(h_cnt >= bagel5_x+28 && h_cnt <= bagel5_x+32 && v_cnt >= bagel5_y+18 && v_cnt <= bagel5_y+20)||(h_cnt >= bagel5_x+4 && h_cnt <= bagel5_x+6 && v_cnt >= bagel5_y+18 && v_cnt <= bagel5_y+20)||(h_cnt >= bagel5_x+6 && h_cnt <= bagel5_x+10 && v_cnt >= bagel5_y+20 && v_cnt <= bagel5_y+22)||(h_cnt >= bagel5_x+12 && h_cnt <= bagel5_x+16 && v_cnt >= bagel5_y+20 && v_cnt <= bagel5_y+22)||(h_cnt >= bagel5_x+26 && h_cnt <= bagel5_x+30 && v_cnt >= bagel5_y+20 && v_cnt <= bagel5_y+22)||(h_cnt >= bagel5_x+34 && h_cnt <= bagel5_x+36 && v_cnt >= bagel5_y+20 && v_cnt <= bagel5_y+22)||(h_cnt >= bagel5_x+4 && h_cnt <= bagel5_x+6 && v_cnt >= bagel5_y+22 && v_cnt <= bagel5_y+24)||(h_cnt >= bagel5_x+8 && h_cnt <= bagel5_x+12 && v_cnt >= bagel5_y+22 && v_cnt <= bagel5_y+24)||(h_cnt >= bagel5_x+14 && h_cnt <= bagel5_x+22 && v_cnt >= bagel5_y+22 && v_cnt <= bagel5_y+24)||(h_cnt >= bagel5_x+24 && h_cnt <= bagel5_x+28 && v_cnt >= bagel5_y+22 && v_cnt <= bagel5_y+24)||(h_cnt >= bagel5_x+32 && h_cnt <= bagel5_x+34 && v_cnt >= bagel5_y+22 && v_cnt <= bagel5_y+24)||(h_cnt >= bagel5_x+6 && h_cnt <= bagel5_x+8 && v_cnt >= bagel5_y+24 && v_cnt <= bagel5_y+26)||(h_cnt >= bagel5_x+12 && h_cnt <= bagel5_x+24 && v_cnt >= bagel5_y+24 && v_cnt <= bagel5_y+26)||(h_cnt >= bagel5_x+30 && h_cnt <= bagel5_x+32 && v_cnt >= bagel5_y+24 && v_cnt <= bagel5_y+26)||(h_cnt >= bagel5_x+8 && h_cnt <= bagel5_x+10 && v_cnt >= bagel5_y+26 && v_cnt <= bagel5_y+28)||(h_cnt >= bagel5_x+28 && h_cnt <= bagel5_x+30 && v_cnt >= bagel5_y+26 && v_cnt <= bagel5_y+28)||(h_cnt >= bagel5_x+12 && h_cnt <= bagel5_x+14 && v_cnt >= bagel5_y+28 && v_cnt <= bagel5_y+30)||(h_cnt >= bagel5_x+24 && h_cnt <= bagel5_x+26 && v_cnt >= bagel5_y+28 && v_cnt <= bagel5_y+30))
					{vgaRed, vgaGreen, vgaBlue} = 12'hf9c; // baby pink
				else if((h_cnt >= bagel5_x+16 && h_cnt <= bagel5_x+24 && v_cnt >= bagel5_y+2 && v_cnt <= bagel5_y+4)||(h_cnt >= bagel5_x+10 && h_cnt <= bagel5_x+26 && v_cnt >= bagel5_y+4 && v_cnt <= bagel5_y+6)||(h_cnt >= bagel5_x+8 && h_cnt <= bagel5_x+14 && v_cnt >= bagel5_y+6 && v_cnt <= bagel5_y+8)||(h_cnt >= bagel5_x+26 && h_cnt <= bagel5_x+28 && v_cnt >= bagel5_y+6 && v_cnt <= bagel5_y+20)||(h_cnt >= bagel5_x+28 && h_cnt <= bagel5_x+30 && v_cnt >= bagel5_y+10 && v_cnt <= bagel5_y+18)||(h_cnt >= bagel5_x+24 && h_cnt <= bagel5_x+26 && v_cnt >= bagel5_y+14 && v_cnt <= bagel5_y+22)||(h_cnt >= bagel5_x+14 && h_cnt <= bagel5_x+24 && v_cnt >= bagel5_y+10 && v_cnt <= bagel5_y+14)||(h_cnt >= bagel5_x+4 && h_cnt <= bagel5_x+10 && v_cnt >= bagel5_y+10 && v_cnt <= bagel5_y+18)||(h_cnt >= bagel5_x+2 && h_cnt <= bagel5_x+4 && v_cnt >= bagel5_y+12 && v_cnt <= bagel5_y+24)||(h_cnt >= bagel5_x+6 && h_cnt <= bagel5_x+10 && v_cnt >= bagel5_y+18 && v_cnt <= bagel5_y+20)||(h_cnt >= bagel5_x+4 && h_cnt <= bagel5_x+6 && v_cnt >= bagel5_y+20 && v_cnt <= bagel5_y+22)||(h_cnt >= bagel5_x+34 && h_cnt <= bagel5_x+36 && v_cnt >= bagel5_y+12 && v_cnt <= bagel5_y+20)||(h_cnt >= bagel5_x+22 && h_cnt <= bagel5_x+24 && v_cnt >= bagel5_y+14 && v_cnt <= bagel5_y+16)||(h_cnt >= bagel5_x+14 && h_cnt <= bagel5_x+18 && v_cnt >= bagel5_y+14 && v_cnt <= bagel5_y+16)||(h_cnt >= bagel5_x+14 && h_cnt <= bagel5_x+16 && v_cnt >= bagel5_y+16 && v_cnt <= bagel5_y+20)||(h_cnt >= bagel5_x+32 && h_cnt <= bagel5_x+34 && v_cnt >= bagel5_y+18 && v_cnt <= bagel5_y+22)||(h_cnt >= bagel5_x+30 && h_cnt <= bagel5_x+32 && v_cnt >= bagel5_y+20 && v_cnt <= bagel5_y+24)||(h_cnt >= bagel5_x+28 && h_cnt <= bagel5_x+30 && v_cnt >= bagel5_y+22 && v_cnt <= bagel5_y+26)||(h_cnt >= bagel5_x+24 && h_cnt <= bagel5_x+28 && v_cnt >= bagel5_y+24 && v_cnt <= bagel5_y+28)||(h_cnt >= bagel5_x+14 && h_cnt <= bagel5_x+26 && v_cnt >= bagel5_y+26 && v_cnt <= bagel5_y+30)||(h_cnt >= bagel5_x+10 && h_cnt <= bagel5_x+14 && v_cnt >= bagel5_y+26 && v_cnt <= bagel5_y+28)||(h_cnt >= bagel5_x+8 && h_cnt <= bagel5_x+12 && v_cnt >= bagel5_y+24 && v_cnt <= bagel5_y+26)||(h_cnt >= bagel5_x+6 && h_cnt <= bagel5_x+12 && v_cnt >= bagel5_y+8 && v_cnt <= bagel5_y+10))
					{vgaRed, vgaGreen, vgaBlue} = 12'hf69; // light pink
				else if((h_cnt >= bagel5_x+12 && h_cnt <= bagel5_x+14 && v_cnt >= bagel5_y+2 && v_cnt <= bagel5_y+4)||(h_cnt >= bagel5_x+28 && h_cnt <= bagel5_x+30 && v_cnt >= bagel5_y+4 && v_cnt <= bagel5_y+6)||(h_cnt >= bagel5_x+30 && h_cnt <= bagel5_x+32 && v_cnt >= bagel5_y+6 && v_cnt <= bagel5_y+8)||(h_cnt >= bagel5_x+32 && h_cnt <= bagel5_x+34 && v_cnt >= bagel5_y+8 && v_cnt <= bagel5_y+10)||(h_cnt >= bagel5_x+10 && h_cnt <= bagel5_x+12 && v_cnt >= bagel5_y+20 && v_cnt <= bagel5_y+22)||(h_cnt >= bagel5_x+16 && h_cnt <= bagel5_x+18 && v_cnt >= bagel5_y+20 && v_cnt <= bagel5_y+22)||(h_cnt >= bagel5_x+22 && h_cnt <= bagel5_x+24 && v_cnt >= bagel5_y+20 && v_cnt <= bagel5_y+24)||(h_cnt >= bagel5_x+6 && h_cnt <= bagel5_x+8 && v_cnt >= bagel5_y+22 && v_cnt <= bagel5_y+24)||(h_cnt >= bagel5_x+32 && h_cnt <= bagel5_x+34 && v_cnt >= bagel5_y+24 && v_cnt <= bagel5_y+28)||(h_cnt >= bagel5_x+34 && h_cnt <= bagel5_x+36 && v_cnt >= bagel5_y+22 && v_cnt <= bagel5_y+24))
					{vgaRed, vgaGreen, vgaBlue} = 12'hf48; // dark pink
				else if((h_cnt >= bagel5_x+4 && h_cnt <= bagel5_x+6 && v_cnt >= bagel5_y+24 && v_cnt <= bagel5_y+28)||(h_cnt >= bagel5_x+6 && h_cnt <= bagel5_x+8 && v_cnt >= bagel5_y+26 && v_cnt <= bagel5_y+30)||(h_cnt >= bagel5_x+8 && h_cnt <= bagel5_x+12 && v_cnt >= bagel5_y+28 && v_cnt <= bagel5_y+32)||(h_cnt >= bagel5_x+12 && h_cnt <= bagel5_x+26 && v_cnt >= bagel5_y+30 && v_cnt <= bagel5_y+34)||(h_cnt >= bagel5_x+26 && h_cnt <= bagel5_x+30 && v_cnt >= bagel5_y+28 && v_cnt <= bagel5_y+32)||(h_cnt >= bagel5_x+30 && h_cnt <= bagel5_x+32 && v_cnt >= bagel5_y+26 && v_cnt <= bagel5_y+30)||(h_cnt >= bagel5_x+4 && h_cnt <= bagel5_x+6 && v_cnt >= bagel5_y+24 && v_cnt <= bagel5_y+28)||(h_cnt >= bagel5_x+12 && h_cnt <= bagel5_x+14 && v_cnt >= bagel5_y+22 && v_cnt <= bagel5_y+24))
					{vgaRed, vgaGreen, vgaBlue} = 12'hfd5; // yellowelse */
				else
					{vgaRed, vgaGreen, vgaBlue} = pixel;
			end
			default:begin
				if(!valid)
					 {vgaRed, vgaGreen, vgaBlue} = 12'h0;
				else
					 {vgaRed, vgaGreen, vgaBlue} = 12'h0;
			end
		endcase
   end   
endmodule
